magic
tech gf180mcuD
magscale 1 10
timestamp 1700882529
<< nwell >>
rect 1258 346880 558742 347744
rect 1258 345312 558742 346176
rect 1258 343744 558742 344608
rect 1258 342176 558742 343040
rect 1258 340608 558742 341472
rect 1258 339040 558742 339904
rect 1258 337472 558742 338336
rect 1258 335904 558742 336768
rect 1258 334336 558742 335200
rect 1258 332768 558742 333632
rect 1258 331200 558742 332064
rect 1258 329632 558742 330496
rect 1258 328064 558742 328928
rect 1258 326496 558742 327360
rect 1258 324928 558742 325792
rect 1258 323360 558742 324224
rect 1258 321792 558742 322656
rect 1258 320224 558742 321088
rect 1258 318656 558742 319520
rect 1258 317088 558742 317952
rect 1258 315520 558742 316384
rect 1258 313952 558742 314816
rect 1258 312384 558742 313248
rect 1258 310816 558742 311680
rect 1258 309248 558742 310112
rect 1258 307680 558742 308544
rect 1258 306112 558742 306976
rect 1258 304544 558742 305408
rect 1258 302976 558742 303840
rect 1258 301408 558742 302272
rect 1258 299840 558742 300704
rect 1258 298272 558742 299136
rect 1258 296704 558742 297568
rect 1258 295136 558742 296000
rect 1258 293568 558742 294432
rect 1258 292000 558742 292864
rect 1258 290432 558742 291296
rect 1258 288864 558742 289728
rect 1258 287296 558742 288160
rect 1258 285728 558742 286592
rect 1258 284160 558742 285024
rect 1258 282592 558742 283456
rect 1258 281024 558742 281888
rect 1258 279456 558742 280320
rect 1258 277888 558742 278752
rect 1258 276320 558742 277184
rect 1258 274752 558742 275616
rect 1258 273184 558742 274048
rect 1258 271616 558742 272480
rect 1258 270048 558742 270912
rect 1258 268480 558742 269344
rect 1258 266912 558742 267776
rect 1258 265344 558742 266208
rect 1258 263776 558742 264640
rect 1258 262208 558742 263072
rect 1258 260640 558742 261504
rect 1258 259072 558742 259936
rect 1258 257504 558742 258368
rect 1258 255936 558742 256800
rect 1258 254368 558742 255232
rect 1258 252800 558742 253664
rect 1258 251232 558742 252096
rect 1258 249664 558742 250528
rect 1258 248096 558742 248960
rect 1258 246528 558742 247392
rect 1258 244960 558742 245824
rect 1258 243392 558742 244256
rect 1258 241824 558742 242688
rect 1258 240256 558742 241120
rect 1258 238688 558742 239552
rect 1258 237120 558742 237984
rect 1258 235552 558742 236416
rect 1258 233984 558742 234848
rect 1258 232416 558742 233280
rect 1258 230848 558742 231712
rect 1258 229280 558742 230144
rect 1258 227712 558742 228576
rect 1258 226144 558742 227008
rect 1258 224576 558742 225440
rect 1258 223008 558742 223872
rect 1258 221440 558742 222304
rect 1258 219872 558742 220736
rect 1258 218304 558742 219168
rect 1258 216736 558742 217600
rect 1258 215168 558742 216032
rect 1258 213600 558742 214464
rect 1258 212032 558742 212896
rect 1258 210464 558742 211328
rect 1258 208896 558742 209760
rect 1258 207328 558742 208192
rect 1258 205760 558742 206624
rect 1258 204192 558742 205056
rect 1258 202624 558742 203488
rect 1258 201056 558742 201920
rect 1258 199488 558742 200352
rect 1258 197920 558742 198784
rect 1258 196352 558742 197216
rect 1258 194784 558742 195648
rect 1258 193216 558742 194080
rect 1258 191648 558742 192512
rect 1258 190080 558742 190944
rect 1258 188512 558742 189376
rect 1258 186944 558742 187808
rect 1258 185376 558742 186240
rect 1258 183808 558742 184672
rect 1258 182240 558742 183104
rect 1258 180672 558742 181536
rect 1258 179104 558742 179968
rect 1258 177536 558742 178400
rect 1258 175968 558742 176832
rect 1258 174400 558742 175264
rect 1258 172832 558742 173696
rect 1258 171264 558742 172128
rect 1258 169696 558742 170560
rect 1258 168128 558742 168992
rect 1258 166560 558742 167424
rect 1258 165831 538728 165856
rect 1258 165017 558742 165831
rect 1258 164992 542984 165017
rect 1258 164263 545302 164288
rect 1258 163449 558742 164263
rect 1258 163424 533869 163449
rect 1258 162695 533240 162720
rect 1258 161881 558742 162695
rect 1258 161856 540094 161881
rect 1258 161127 545224 161152
rect 1258 160313 558742 161127
rect 1258 160288 534429 160313
rect 1258 158745 558742 159584
rect 1258 158720 541261 158745
rect 1258 157991 538013 158016
rect 1258 157177 558742 157991
rect 1258 157152 542381 157177
rect 1258 156423 546887 156448
rect 1258 155584 558742 156423
rect 1258 154855 544397 154880
rect 1258 154041 558742 154855
rect 1258 154016 550936 154041
rect 1258 152448 558742 153312
rect 1258 150880 558742 151744
rect 1258 149312 558742 150176
rect 1258 147744 558742 148608
rect 1258 146176 558742 147040
rect 1258 144608 558742 145472
rect 1258 143040 558742 143904
rect 1258 141472 558742 142336
rect 1258 139904 558742 140768
rect 1258 138336 558742 139200
rect 1258 136768 558742 137632
rect 1258 135200 558742 136064
rect 1258 133632 558742 134496
rect 1258 132064 558742 132928
rect 1258 130496 558742 131360
rect 1258 128928 558742 129792
rect 1258 127360 558742 128224
rect 1258 125792 558742 126656
rect 1258 124224 558742 125088
rect 1258 122656 558742 123520
rect 1258 121088 558742 121952
rect 1258 119520 558742 120384
rect 1258 117952 558742 118816
rect 1258 116384 558742 117248
rect 1258 114816 558742 115680
rect 1258 113248 558742 114112
rect 1258 111680 558742 112544
rect 1258 110112 558742 110976
rect 1258 108544 558742 109408
rect 1258 106976 558742 107840
rect 1258 105408 558742 106272
rect 1258 103840 558742 104704
rect 1258 102272 558742 103136
rect 1258 100704 558742 101568
rect 1258 99136 558742 100000
rect 1258 97568 558742 98432
rect 1258 96000 558742 96864
rect 1258 94432 558742 95296
rect 1258 92864 558742 93728
rect 1258 91296 558742 92160
rect 1258 89728 558742 90592
rect 1258 88160 558742 89024
rect 1258 86592 558742 87456
rect 1258 85024 558742 85888
rect 1258 83456 558742 84320
rect 1258 81888 558742 82752
rect 1258 80320 558742 81184
rect 1258 78752 558742 79616
rect 1258 77184 558742 78048
rect 1258 75616 558742 76480
rect 1258 74048 558742 74912
rect 1258 72480 558742 73344
rect 1258 70912 558742 71776
rect 1258 69344 558742 70208
rect 1258 67776 558742 68640
rect 1258 66208 558742 67072
rect 1258 64640 558742 65504
rect 1258 63072 558742 63936
rect 1258 61504 558742 62368
rect 1258 59936 558742 60800
rect 1258 58368 558742 59232
rect 1258 56800 558742 57664
rect 1258 55232 558742 56096
rect 1258 53664 558742 54528
rect 1258 52096 558742 52960
rect 1258 50528 558742 51392
rect 1258 48960 558742 49824
rect 1258 47392 558742 48256
rect 1258 45824 558742 46688
rect 1258 44256 558742 45120
rect 1258 42688 558742 43552
rect 1258 41120 558742 41984
rect 1258 39552 558742 40416
rect 1258 37984 558742 38848
rect 1258 36416 558742 37280
rect 1258 34848 558742 35712
rect 1258 33280 558742 34144
rect 1258 31712 558742 32576
rect 1258 30144 558742 31008
rect 1258 28576 558742 29440
rect 1258 27008 558742 27872
rect 1258 25440 558742 26304
rect 1258 23872 558742 24736
rect 1258 22304 558742 23168
rect 1258 20736 558742 21600
rect 1258 19168 558742 20032
rect 1258 17600 558742 18464
rect 1258 16032 558742 16896
rect 1258 14464 558742 15328
rect 1258 12896 558742 13760
rect 1258 11328 558742 12192
rect 1258 9760 558742 10624
rect 1258 8192 558742 9056
rect 1258 6624 558742 7488
rect 1258 5056 558742 5920
rect 1258 3488 558742 4352
<< pwell >>
rect 1258 347744 558742 348182
rect 1258 346176 558742 346880
rect 1258 344608 558742 345312
rect 1258 343040 558742 343744
rect 1258 341472 558742 342176
rect 1258 339904 558742 340608
rect 1258 338336 558742 339040
rect 1258 336768 558742 337472
rect 1258 335200 558742 335904
rect 1258 333632 558742 334336
rect 1258 332064 558742 332768
rect 1258 330496 558742 331200
rect 1258 328928 558742 329632
rect 1258 327360 558742 328064
rect 1258 325792 558742 326496
rect 1258 324224 558742 324928
rect 1258 322656 558742 323360
rect 1258 321088 558742 321792
rect 1258 319520 558742 320224
rect 1258 317952 558742 318656
rect 1258 316384 558742 317088
rect 1258 314816 558742 315520
rect 1258 313248 558742 313952
rect 1258 311680 558742 312384
rect 1258 310112 558742 310816
rect 1258 308544 558742 309248
rect 1258 306976 558742 307680
rect 1258 305408 558742 306112
rect 1258 303840 558742 304544
rect 1258 302272 558742 302976
rect 1258 300704 558742 301408
rect 1258 299136 558742 299840
rect 1258 297568 558742 298272
rect 1258 296000 558742 296704
rect 1258 294432 558742 295136
rect 1258 292864 558742 293568
rect 1258 291296 558742 292000
rect 1258 289728 558742 290432
rect 1258 288160 558742 288864
rect 1258 286592 558742 287296
rect 1258 285024 558742 285728
rect 1258 283456 558742 284160
rect 1258 281888 558742 282592
rect 1258 280320 558742 281024
rect 1258 278752 558742 279456
rect 1258 277184 558742 277888
rect 1258 275616 558742 276320
rect 1258 274048 558742 274752
rect 1258 272480 558742 273184
rect 1258 270912 558742 271616
rect 1258 269344 558742 270048
rect 1258 267776 558742 268480
rect 1258 266208 558742 266912
rect 1258 264640 558742 265344
rect 1258 263072 558742 263776
rect 1258 261504 558742 262208
rect 1258 259936 558742 260640
rect 1258 258368 558742 259072
rect 1258 256800 558742 257504
rect 1258 255232 558742 255936
rect 1258 253664 558742 254368
rect 1258 252096 558742 252800
rect 1258 250528 558742 251232
rect 1258 248960 558742 249664
rect 1258 247392 558742 248096
rect 1258 245824 558742 246528
rect 1258 244256 558742 244960
rect 1258 242688 558742 243392
rect 1258 241120 558742 241824
rect 1258 239552 558742 240256
rect 1258 237984 558742 238688
rect 1258 236416 558742 237120
rect 1258 234848 558742 235552
rect 1258 233280 558742 233984
rect 1258 231712 558742 232416
rect 1258 230144 558742 230848
rect 1258 228576 558742 229280
rect 1258 227008 558742 227712
rect 1258 225440 558742 226144
rect 1258 223872 558742 224576
rect 1258 222304 558742 223008
rect 1258 220736 558742 221440
rect 1258 219168 558742 219872
rect 1258 217600 558742 218304
rect 1258 216032 558742 216736
rect 1258 214464 558742 215168
rect 1258 212896 558742 213600
rect 1258 211328 558742 212032
rect 1258 209760 558742 210464
rect 1258 208192 558742 208896
rect 1258 206624 558742 207328
rect 1258 205056 558742 205760
rect 1258 203488 558742 204192
rect 1258 201920 558742 202624
rect 1258 200352 558742 201056
rect 1258 198784 558742 199488
rect 1258 197216 558742 197920
rect 1258 195648 558742 196352
rect 1258 194080 558742 194784
rect 1258 192512 558742 193216
rect 1258 190944 558742 191648
rect 1258 189376 558742 190080
rect 1258 187808 558742 188512
rect 1258 186240 558742 186944
rect 1258 184672 558742 185376
rect 1258 183104 558742 183808
rect 1258 181536 558742 182240
rect 1258 179968 558742 180672
rect 1258 178400 558742 179104
rect 1258 176832 558742 177536
rect 1258 175264 558742 175968
rect 1258 173696 558742 174400
rect 1258 172128 558742 172832
rect 1258 170560 558742 171264
rect 1258 168992 558742 169696
rect 1258 167424 558742 168128
rect 1258 165856 558742 166560
rect 1258 164288 558742 164992
rect 1258 162720 558742 163424
rect 1258 161152 558742 161856
rect 1258 159584 558742 160288
rect 1258 158016 558742 158720
rect 1258 156448 558742 157152
rect 1258 154880 558742 155584
rect 1258 153312 558742 154016
rect 1258 151744 558742 152448
rect 1258 150176 558742 150880
rect 1258 148608 558742 149312
rect 1258 147040 558742 147744
rect 1258 145472 558742 146176
rect 1258 143904 558742 144608
rect 1258 142336 558742 143040
rect 1258 140768 558742 141472
rect 1258 139200 558742 139904
rect 1258 137632 558742 138336
rect 1258 136064 558742 136768
rect 1258 134496 558742 135200
rect 1258 132928 558742 133632
rect 1258 131360 558742 132064
rect 1258 129792 558742 130496
rect 1258 128224 558742 128928
rect 1258 126656 558742 127360
rect 1258 125088 558742 125792
rect 1258 123520 558742 124224
rect 1258 121952 558742 122656
rect 1258 120384 558742 121088
rect 1258 118816 558742 119520
rect 1258 117248 558742 117952
rect 1258 115680 558742 116384
rect 1258 114112 558742 114816
rect 1258 112544 558742 113248
rect 1258 110976 558742 111680
rect 1258 109408 558742 110112
rect 1258 107840 558742 108544
rect 1258 106272 558742 106976
rect 1258 104704 558742 105408
rect 1258 103136 558742 103840
rect 1258 101568 558742 102272
rect 1258 100000 558742 100704
rect 1258 98432 558742 99136
rect 1258 96864 558742 97568
rect 1258 95296 558742 96000
rect 1258 93728 558742 94432
rect 1258 92160 558742 92864
rect 1258 90592 558742 91296
rect 1258 89024 558742 89728
rect 1258 87456 558742 88160
rect 1258 85888 558742 86592
rect 1258 84320 558742 85024
rect 1258 82752 558742 83456
rect 1258 81184 558742 81888
rect 1258 79616 558742 80320
rect 1258 78048 558742 78752
rect 1258 76480 558742 77184
rect 1258 74912 558742 75616
rect 1258 73344 558742 74048
rect 1258 71776 558742 72480
rect 1258 70208 558742 70912
rect 1258 68640 558742 69344
rect 1258 67072 558742 67776
rect 1258 65504 558742 66208
rect 1258 63936 558742 64640
rect 1258 62368 558742 63072
rect 1258 60800 558742 61504
rect 1258 59232 558742 59936
rect 1258 57664 558742 58368
rect 1258 56096 558742 56800
rect 1258 54528 558742 55232
rect 1258 52960 558742 53664
rect 1258 51392 558742 52096
rect 1258 49824 558742 50528
rect 1258 48256 558742 48960
rect 1258 46688 558742 47392
rect 1258 45120 558742 45824
rect 1258 43552 558742 44256
rect 1258 41984 558742 42688
rect 1258 40416 558742 41120
rect 1258 38848 558742 39552
rect 1258 37280 558742 37984
rect 1258 35712 558742 36416
rect 1258 34144 558742 34848
rect 1258 32576 558742 33280
rect 1258 31008 558742 31712
rect 1258 29440 558742 30144
rect 1258 27872 558742 28576
rect 1258 26304 558742 27008
rect 1258 24736 558742 25440
rect 1258 23168 558742 23872
rect 1258 21600 558742 22304
rect 1258 20032 558742 20736
rect 1258 18464 558742 19168
rect 1258 16896 558742 17600
rect 1258 15328 558742 16032
rect 1258 13760 558742 14464
rect 1258 12192 558742 12896
rect 1258 10624 558742 11328
rect 1258 9056 558742 9760
rect 1258 7488 558742 8192
rect 1258 5920 558742 6624
rect 1258 4352 558742 5056
rect 1258 3050 558742 3488
<< obsm1 >>
rect 1344 3076 558656 348156
<< metal2 >>
rect 139776 0 139888 800
rect 419776 0 419888 800
<< obsm2 >>
rect 4476 860 558292 348134
rect 4476 800 139716 860
rect 139948 800 419716 860
rect 419948 800 558292 860
<< metal3 >>
rect 559200 326368 560000 326480
rect 559200 276192 560000 276304
rect 559200 226016 560000 226128
rect 559200 175840 560000 175952
rect 559200 125664 560000 125776
rect 559200 75488 560000 75600
rect 559200 25312 560000 25424
<< obsm3 >>
rect 4466 326540 559200 348124
rect 4466 326308 559140 326540
rect 4466 276364 559200 326308
rect 4466 276132 559140 276364
rect 4466 226188 559200 276132
rect 4466 225956 559140 226188
rect 4466 176012 559200 225956
rect 4466 175780 559140 176012
rect 4466 125836 559200 175780
rect 4466 125604 559140 125836
rect 4466 75660 559200 125604
rect 4466 75428 559140 75660
rect 4466 25484 559200 75428
rect 4466 25252 559140 25484
rect 4466 3108 559200 25252
<< metal4 >>
rect 4448 3076 4768 348156
rect 19808 3076 20128 348156
rect 35168 3076 35488 348156
rect 50528 3076 50848 348156
rect 65888 3076 66208 348156
rect 81248 3076 81568 348156
rect 96608 3076 96928 348156
rect 111968 3076 112288 348156
rect 127328 3076 127648 348156
rect 142688 3076 143008 348156
rect 158048 3076 158368 348156
rect 173408 3076 173728 348156
rect 188768 3076 189088 348156
rect 204128 3076 204448 348156
rect 219488 3076 219808 348156
rect 234848 3076 235168 348156
rect 250208 3076 250528 348156
rect 265568 3076 265888 348156
rect 280928 3076 281248 348156
rect 296288 3076 296608 348156
rect 311648 3076 311968 348156
rect 327008 3076 327328 348156
rect 342368 3076 342688 348156
rect 357728 3076 358048 348156
rect 373088 3076 373408 348156
rect 388448 3076 388768 348156
rect 403808 3076 404128 348156
rect 419168 3076 419488 348156
rect 434528 3076 434848 348156
rect 449888 3076 450208 348156
rect 465248 3076 465568 348156
rect 480608 3076 480928 348156
rect 495968 3076 496288 348156
rect 511328 3076 511648 348156
rect 526688 3076 527008 348156
rect 542048 3076 542368 348156
rect 557408 3076 557728 348156
<< obsm4 >>
rect 548940 155922 548996 156894
<< labels >>
rlabel metal3 s 559200 326368 560000 326480 6 clk_fin
port 1 nsew signal input
rlabel metal3 s 559200 226016 560000 226128 6 freq_select[0]
port 2 nsew signal input
rlabel metal3 s 559200 276192 560000 276304 6 freq_select[1]
port 3 nsew signal input
rlabel metal3 s 559200 25312 560000 25424 6 io_oeb[0]
port 4 nsew signal output
rlabel metal3 s 559200 125664 560000 125776 6 io_oeb[1]
port 5 nsew signal output
rlabel metal3 s 559200 75488 560000 75600 6 io_out[0]
port 6 nsew signal output
rlabel metal3 s 559200 175840 560000 175952 6 io_out[1]
port 7 nsew signal output
rlabel metal4 s 4448 3076 4768 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 526688 3076 527008 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 557408 3076 557728 348156 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 542048 3076 542368 348156 6 vss
port 9 nsew ground bidirectional
rlabel metal2 s 139776 0 139888 800 6 wb_clk_i
port 10 nsew signal input
rlabel metal2 s 419776 0 419888 800 6 wb_rst_i
port 11 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15130466
string GDS_FILE /home/oe23ranan/dpll-project/openlane/dpll/runs/23_11_25_12_17/results/signoff/dpll.magic.gds
string GDS_START 185340
<< end >>

