VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO anan_logo
  CLASS BLOCK ;
  FOREIGN anan_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 352.200 ;
  PIN vdd
    PORT
      LAYER Metal5 ;
        RECT 147.500 342.600 152.500 344.700 ;
        RECT 125.000 342.000 175.000 342.600 ;
        RECT 124.800 341.400 175.200 342.000 ;
        RECT 124.600 340.800 175.400 341.400 ;
        RECT 124.300 340.200 175.700 340.800 ;
        RECT 124.100 339.600 175.900 340.200 ;
        RECT 123.900 339.000 176.100 339.600 ;
        RECT 123.600 338.400 176.400 339.000 ;
        RECT 123.400 337.800 176.600 338.400 ;
        RECT 123.200 337.200 176.800 337.800 ;
        RECT 123.000 336.600 177.000 337.200 ;
        RECT 122.800 336.000 177.200 336.600 ;
        RECT 122.500 335.400 177.500 336.000 ;
        RECT 122.300 334.800 177.700 335.400 ;
        RECT 122.100 334.200 177.900 334.800 ;
        RECT 121.800 333.600 178.200 334.200 ;
        RECT 121.600 333.000 178.400 333.600 ;
        RECT 121.400 332.400 178.600 333.000 ;
        RECT 121.200 331.800 178.800 332.400 ;
        RECT 120.900 331.200 179.000 331.800 ;
        RECT 120.700 330.600 179.300 331.200 ;
        RECT 120.500 330.000 179.500 330.600 ;
        RECT 120.300 329.400 179.700 330.000 ;
        RECT 120.100 328.800 180.000 329.400 ;
        RECT 119.800 328.200 180.200 328.800 ;
        RECT 119.600 327.600 180.400 328.200 ;
        RECT 119.400 327.000 180.600 327.600 ;
        RECT 119.200 326.400 180.800 327.000 ;
        RECT 118.900 325.800 181.100 326.400 ;
        RECT 118.700 325.200 181.300 325.800 ;
        RECT 118.500 324.600 181.500 325.200 ;
        RECT 118.200 324.000 181.800 324.600 ;
        RECT 118.000 323.400 182.000 324.000 ;
        RECT 117.800 322.800 182.200 323.400 ;
        RECT 117.600 322.200 182.400 322.800 ;
        RECT 117.400 321.600 182.600 322.200 ;
        RECT 117.100 321.000 182.900 321.600 ;
        RECT 116.900 320.400 183.100 321.000 ;
        RECT 116.700 319.800 183.300 320.400 ;
        RECT 116.400 319.200 183.600 319.800 ;
        RECT 116.200 318.600 183.800 319.200 ;
        RECT 116.000 318.000 184.000 318.600 ;
        RECT 115.800 317.400 184.200 318.000 ;
        RECT 115.600 316.800 184.400 317.400 ;
        RECT 115.300 316.200 184.700 316.800 ;
        RECT 115.100 315.600 184.900 316.200 ;
        RECT 114.900 315.000 185.100 315.600 ;
        RECT 114.600 314.400 185.400 315.000 ;
        RECT 114.400 313.800 185.600 314.400 ;
        RECT 114.200 313.200 185.800 313.800 ;
        RECT 114.000 312.600 186.000 313.200 ;
        RECT 113.800 312.000 186.200 312.600 ;
        RECT 113.500 311.400 186.500 312.000 ;
        RECT 113.300 310.800 186.700 311.400 ;
        RECT 113.100 310.200 186.900 310.800 ;
        RECT 112.800 309.600 187.200 310.200 ;
        RECT 112.600 309.000 187.400 309.600 ;
        RECT 112.400 308.400 187.600 309.000 ;
        RECT 112.200 307.800 187.800 308.400 ;
        RECT 111.900 307.200 188.000 307.800 ;
        RECT 111.700 306.600 188.300 307.200 ;
        RECT 111.500 306.000 188.500 306.600 ;
        RECT 111.300 305.400 188.700 306.000 ;
        RECT 111.100 304.800 189.000 305.400 ;
        RECT 110.800 304.200 189.200 304.800 ;
        RECT 110.600 303.600 189.400 304.200 ;
        RECT 110.400 303.000 189.600 303.600 ;
        RECT 110.200 302.400 189.800 303.000 ;
        RECT 109.900 301.800 190.100 302.400 ;
        RECT 109.700 301.200 190.300 301.800 ;
        RECT 109.500 300.600 190.500 301.200 ;
        RECT 109.200 300.000 190.800 300.600 ;
        RECT 109.000 299.400 191.000 300.000 ;
        RECT 108.800 298.800 191.200 299.400 ;
        RECT 108.600 298.200 191.400 298.800 ;
        RECT 108.400 297.600 191.600 298.200 ;
        RECT 108.100 297.000 191.900 297.600 ;
        RECT 107.900 296.400 192.100 297.000 ;
        RECT 107.700 295.800 192.300 296.400 ;
        RECT 107.400 295.200 192.600 295.800 ;
        RECT 107.200 294.600 192.800 295.200 ;
        RECT 107.000 294.000 193.000 294.600 ;
        RECT 106.800 293.400 193.200 294.000 ;
        RECT 106.600 292.800 193.400 293.400 ;
        RECT 106.300 292.200 193.700 292.800 ;
        RECT 106.100 291.600 193.900 292.200 ;
        RECT 105.900 291.000 194.100 291.600 ;
        RECT 105.600 290.400 194.400 291.000 ;
        RECT 105.400 289.800 194.600 290.400 ;
        RECT 105.200 289.200 194.800 289.800 ;
        RECT 105.000 288.600 195.000 289.200 ;
        RECT 104.800 288.000 195.200 288.600 ;
        RECT 104.500 287.400 195.500 288.000 ;
        RECT 104.300 286.800 195.700 287.400 ;
        RECT 104.100 286.200 195.900 286.800 ;
        RECT 103.800 285.600 196.200 286.200 ;
        RECT 103.600 285.000 196.400 285.600 ;
        RECT 103.400 284.400 196.600 285.000 ;
        RECT 103.200 283.800 196.800 284.400 ;
        RECT 103.000 283.200 197.000 283.800 ;
        RECT 102.700 282.600 197.300 283.200 ;
        RECT 102.500 282.000 197.500 282.600 ;
        RECT 102.300 281.400 197.700 282.000 ;
        RECT 102.000 280.800 198.000 281.400 ;
        RECT 101.800 280.200 198.200 280.800 ;
        RECT 101.600 279.600 198.400 280.200 ;
        RECT 101.400 279.000 198.600 279.600 ;
        RECT 101.200 278.400 198.800 279.000 ;
        RECT 100.900 277.800 199.100 278.400 ;
        RECT 100.700 277.200 199.300 277.800 ;
        RECT 100.500 276.600 199.500 277.200 ;
        RECT 100.200 276.000 199.800 276.600 ;
        RECT 100.000 275.400 200.000 276.000 ;
        RECT 99.800 275.200 200.200 275.400 ;
        RECT 99.800 274.800 149.800 275.200 ;
        RECT 99.600 274.600 149.800 274.800 ;
        RECT 150.200 274.800 200.200 275.200 ;
        RECT 150.200 274.600 200.400 274.800 ;
        RECT 99.600 274.200 149.600 274.600 ;
        RECT 99.400 274.000 149.600 274.200 ;
        RECT 150.400 274.200 200.400 274.600 ;
        RECT 150.400 274.000 200.600 274.200 ;
        RECT 99.400 273.600 149.400 274.000 ;
        RECT 99.100 273.400 149.400 273.600 ;
        RECT 150.600 273.600 200.600 274.000 ;
        RECT 150.600 273.400 200.900 273.600 ;
        RECT 99.100 273.000 149.100 273.400 ;
        RECT 98.900 272.800 149.100 273.000 ;
        RECT 150.900 273.000 200.900 273.400 ;
        RECT 150.900 272.800 201.100 273.000 ;
        RECT 98.900 272.400 148.900 272.800 ;
        RECT 98.700 272.200 148.900 272.400 ;
        RECT 151.100 272.400 201.100 272.800 ;
        RECT 151.100 272.200 201.300 272.400 ;
        RECT 98.700 271.800 148.700 272.200 ;
        RECT 98.400 271.600 148.700 271.800 ;
        RECT 151.300 271.800 201.300 272.200 ;
        RECT 151.300 271.600 201.600 271.800 ;
        RECT 98.400 271.200 148.400 271.600 ;
        RECT 98.200 271.000 148.400 271.200 ;
        RECT 151.600 271.200 201.600 271.600 ;
        RECT 151.600 271.000 201.800 271.200 ;
        RECT 98.200 270.600 148.200 271.000 ;
        RECT 98.000 270.400 148.200 270.600 ;
        RECT 151.800 270.600 201.800 271.000 ;
        RECT 151.800 270.400 202.000 270.600 ;
        RECT 98.000 270.000 148.000 270.400 ;
        RECT 97.800 269.800 148.000 270.000 ;
        RECT 152.000 270.000 202.000 270.400 ;
        RECT 152.000 269.800 202.200 270.000 ;
        RECT 97.800 269.400 147.800 269.800 ;
        RECT 97.600 269.200 147.800 269.400 ;
        RECT 152.200 269.400 202.200 269.800 ;
        RECT 152.200 269.200 202.400 269.400 ;
        RECT 97.600 268.800 147.600 269.200 ;
        RECT 97.300 268.600 147.600 268.800 ;
        RECT 152.400 268.800 202.400 269.200 ;
        RECT 152.400 268.600 202.700 268.800 ;
        RECT 97.300 268.200 147.300 268.600 ;
        RECT 97.100 268.000 147.300 268.200 ;
        RECT 152.700 268.200 202.700 268.600 ;
        RECT 152.700 268.000 202.900 268.200 ;
        RECT 97.100 267.600 147.100 268.000 ;
        RECT 96.900 267.400 147.100 267.600 ;
        RECT 152.900 267.600 202.900 268.000 ;
        RECT 152.900 267.400 203.100 267.600 ;
        RECT 96.900 267.000 146.900 267.400 ;
        RECT 96.600 266.800 146.900 267.000 ;
        RECT 153.100 267.000 203.100 267.400 ;
        RECT 153.100 266.800 203.400 267.000 ;
        RECT 96.600 266.400 146.600 266.800 ;
        RECT 96.400 266.200 146.600 266.400 ;
        RECT 153.400 266.400 203.400 266.800 ;
        RECT 153.400 266.200 203.600 266.400 ;
        RECT 96.400 265.800 146.400 266.200 ;
        RECT 96.200 265.600 146.400 265.800 ;
        RECT 153.600 265.800 203.600 266.200 ;
        RECT 153.600 265.600 203.800 265.800 ;
        RECT 96.200 265.200 146.200 265.600 ;
        RECT 96.000 265.000 146.200 265.200 ;
        RECT 153.800 265.200 203.800 265.600 ;
        RECT 153.800 265.000 204.000 265.200 ;
        RECT 96.000 264.600 146.000 265.000 ;
        RECT 95.800 264.400 146.000 264.600 ;
        RECT 154.000 264.600 204.000 265.000 ;
        RECT 154.000 264.400 204.200 264.600 ;
        RECT 95.800 264.000 145.800 264.400 ;
        RECT 95.500 263.800 145.800 264.000 ;
        RECT 154.200 264.000 204.200 264.400 ;
        RECT 154.200 263.800 204.500 264.000 ;
        RECT 95.500 263.400 145.500 263.800 ;
        RECT 95.300 263.200 145.500 263.400 ;
        RECT 154.500 263.400 204.500 263.800 ;
        RECT 154.500 263.200 204.700 263.400 ;
        RECT 95.300 262.800 145.300 263.200 ;
        RECT 95.100 262.600 145.300 262.800 ;
        RECT 154.700 262.800 204.700 263.200 ;
        RECT 154.700 262.600 204.900 262.800 ;
        RECT 95.100 262.200 145.100 262.600 ;
        RECT 94.800 262.000 145.100 262.200 ;
        RECT 154.900 262.200 204.900 262.600 ;
        RECT 154.900 262.000 205.200 262.200 ;
        RECT 94.800 261.600 144.800 262.000 ;
        RECT 94.600 261.400 144.800 261.600 ;
        RECT 155.200 261.600 205.200 262.000 ;
        RECT 155.200 261.400 205.400 261.600 ;
        RECT 94.600 261.000 144.600 261.400 ;
        RECT 94.400 260.800 144.600 261.000 ;
        RECT 155.400 261.000 205.400 261.400 ;
        RECT 155.400 260.800 205.600 261.000 ;
        RECT 94.400 260.400 144.400 260.800 ;
        RECT 94.200 260.200 144.400 260.400 ;
        RECT 155.600 260.400 205.600 260.800 ;
        RECT 155.600 260.200 205.800 260.400 ;
        RECT 94.200 259.800 144.200 260.200 ;
        RECT 94.000 259.600 144.200 259.800 ;
        RECT 155.800 259.800 205.800 260.200 ;
        RECT 155.800 259.600 206.000 259.800 ;
        RECT 94.000 259.200 144.000 259.600 ;
        RECT 93.700 259.000 144.000 259.200 ;
        RECT 156.000 259.200 206.000 259.600 ;
        RECT 156.000 259.000 206.300 259.200 ;
        RECT 93.700 258.600 143.700 259.000 ;
        RECT 93.500 258.400 143.700 258.600 ;
        RECT 156.300 258.600 206.300 259.000 ;
        RECT 156.300 258.400 206.500 258.600 ;
        RECT 93.500 258.000 143.500 258.400 ;
        RECT 93.300 257.800 143.500 258.000 ;
        RECT 156.500 258.000 206.500 258.400 ;
        RECT 156.500 257.800 206.700 258.000 ;
        RECT 93.300 257.400 143.300 257.800 ;
        RECT 93.000 257.200 143.300 257.400 ;
        RECT 156.700 257.400 206.700 257.800 ;
        RECT 156.700 257.200 207.000 257.400 ;
        RECT 93.000 256.800 143.000 257.200 ;
        RECT 92.800 256.600 143.000 256.800 ;
        RECT 157.000 256.800 207.000 257.200 ;
        RECT 157.000 256.600 207.200 256.800 ;
        RECT 92.800 256.200 142.800 256.600 ;
        RECT 92.600 256.000 142.800 256.200 ;
        RECT 157.200 256.200 207.200 256.600 ;
        RECT 157.200 256.000 207.400 256.200 ;
        RECT 92.600 255.600 142.600 256.000 ;
        RECT 92.400 255.400 142.600 255.600 ;
        RECT 157.400 255.600 207.400 256.000 ;
        RECT 157.400 255.400 207.600 255.600 ;
        RECT 92.400 255.000 142.400 255.400 ;
        RECT 92.200 254.800 142.400 255.000 ;
        RECT 157.600 255.000 207.600 255.400 ;
        RECT 157.600 254.800 207.800 255.000 ;
        RECT 92.200 254.400 142.200 254.800 ;
        RECT 91.900 254.200 142.200 254.400 ;
        RECT 157.800 254.400 207.800 254.800 ;
        RECT 157.800 254.200 208.100 254.400 ;
        RECT 91.900 253.800 141.900 254.200 ;
        RECT 91.700 253.600 141.900 253.800 ;
        RECT 158.100 253.800 208.100 254.200 ;
        RECT 158.100 253.600 208.300 253.800 ;
        RECT 91.700 253.200 141.700 253.600 ;
        RECT 91.500 253.000 141.700 253.200 ;
        RECT 158.300 253.200 208.300 253.600 ;
        RECT 158.300 253.000 208.500 253.200 ;
        RECT 91.500 252.600 141.500 253.000 ;
        RECT 91.200 252.400 141.500 252.600 ;
        RECT 158.500 252.600 208.500 253.000 ;
        RECT 158.500 252.400 208.800 252.600 ;
        RECT 91.200 252.000 141.200 252.400 ;
        RECT 91.000 251.800 141.200 252.000 ;
        RECT 158.800 252.000 208.800 252.400 ;
        RECT 158.800 251.800 209.000 252.000 ;
        RECT 91.000 251.400 141.000 251.800 ;
        RECT 90.800 251.200 141.000 251.400 ;
        RECT 159.000 251.400 209.000 251.800 ;
        RECT 159.000 251.200 209.200 251.400 ;
        RECT 90.800 250.800 140.800 251.200 ;
        RECT 90.600 250.600 140.800 250.800 ;
        RECT 159.200 250.800 209.200 251.200 ;
        RECT 159.200 250.600 209.400 250.800 ;
        RECT 90.600 250.200 140.600 250.600 ;
        RECT 90.400 250.000 140.600 250.200 ;
        RECT 159.400 250.200 209.400 250.600 ;
        RECT 159.400 250.000 209.600 250.200 ;
        RECT 90.400 249.600 140.400 250.000 ;
        RECT 90.100 249.400 140.400 249.600 ;
        RECT 159.600 249.600 209.600 250.000 ;
        RECT 159.600 249.400 209.900 249.600 ;
        RECT 90.100 249.000 140.100 249.400 ;
        RECT 89.900 248.800 140.100 249.000 ;
        RECT 159.900 249.000 209.900 249.400 ;
        RECT 159.900 248.800 210.100 249.000 ;
        RECT 89.900 248.400 139.900 248.800 ;
        RECT 89.700 248.200 139.900 248.400 ;
        RECT 160.100 248.400 210.100 248.800 ;
        RECT 160.100 248.200 210.300 248.400 ;
        RECT 89.700 247.800 139.700 248.200 ;
        RECT 89.400 247.600 139.700 247.800 ;
        RECT 160.300 247.800 210.300 248.200 ;
        RECT 160.300 247.600 210.600 247.800 ;
        RECT 89.400 247.200 139.400 247.600 ;
        RECT 89.200 247.000 139.400 247.200 ;
        RECT 160.600 247.200 210.600 247.600 ;
        RECT 160.600 247.000 210.800 247.200 ;
        RECT 89.200 246.600 139.200 247.000 ;
        RECT 89.000 246.400 139.200 246.600 ;
        RECT 160.800 246.600 210.800 247.000 ;
        RECT 160.800 246.400 211.000 246.600 ;
        RECT 89.000 246.000 139.000 246.400 ;
        RECT 88.800 245.800 139.000 246.000 ;
        RECT 161.000 246.000 211.000 246.400 ;
        RECT 161.000 245.800 211.200 246.000 ;
        RECT 88.800 245.400 138.800 245.800 ;
        RECT 88.600 245.200 138.800 245.400 ;
        RECT 161.200 245.400 211.200 245.800 ;
        RECT 161.200 245.200 211.400 245.400 ;
        RECT 88.600 244.800 138.600 245.200 ;
        RECT 88.300 244.600 138.600 244.800 ;
        RECT 161.400 244.800 211.400 245.200 ;
        RECT 161.400 244.600 211.700 244.800 ;
        RECT 88.300 244.200 138.300 244.600 ;
        RECT 88.100 244.000 138.300 244.200 ;
        RECT 161.700 244.200 211.700 244.600 ;
        RECT 161.700 244.000 211.900 244.200 ;
        RECT 88.100 243.600 138.100 244.000 ;
        RECT 87.900 243.400 138.100 243.600 ;
        RECT 161.900 243.600 211.900 244.000 ;
        RECT 161.900 243.400 212.100 243.600 ;
        RECT 87.900 243.000 137.900 243.400 ;
        RECT 87.600 242.800 137.900 243.000 ;
        RECT 162.100 243.000 212.100 243.400 ;
        RECT 162.100 242.800 212.400 243.000 ;
        RECT 87.600 242.400 137.600 242.800 ;
        RECT 87.400 242.200 137.600 242.400 ;
        RECT 162.400 242.400 212.400 242.800 ;
        RECT 162.400 242.200 212.600 242.400 ;
        RECT 87.400 241.800 137.400 242.200 ;
        RECT 87.200 241.600 137.400 241.800 ;
        RECT 162.600 241.800 212.600 242.200 ;
        RECT 162.600 241.600 212.800 241.800 ;
        RECT 87.200 241.200 137.200 241.600 ;
        RECT 87.000 241.000 137.200 241.200 ;
        RECT 162.800 241.200 212.800 241.600 ;
        RECT 162.800 241.000 213.000 241.200 ;
        RECT 87.000 240.600 137.000 241.000 ;
        RECT 86.800 240.400 137.000 240.600 ;
        RECT 163.000 240.600 213.000 241.000 ;
        RECT 163.000 240.400 213.200 240.600 ;
        RECT 86.800 240.000 136.800 240.400 ;
        RECT 86.500 239.800 136.800 240.000 ;
        RECT 163.200 240.000 213.200 240.400 ;
        RECT 163.200 239.800 213.500 240.000 ;
        RECT 86.500 239.400 136.500 239.800 ;
        RECT 86.300 239.200 136.500 239.400 ;
        RECT 163.500 239.400 213.500 239.800 ;
        RECT 163.500 239.200 213.700 239.400 ;
        RECT 86.300 238.800 136.300 239.200 ;
        RECT 86.100 238.600 136.300 238.800 ;
        RECT 163.700 238.800 213.700 239.200 ;
        RECT 163.700 238.600 213.900 238.800 ;
        RECT 86.100 238.200 136.100 238.600 ;
        RECT 85.800 238.000 136.100 238.200 ;
        RECT 163.900 238.200 213.900 238.600 ;
        RECT 163.900 238.000 214.200 238.200 ;
        RECT 85.800 237.600 135.800 238.000 ;
        RECT 85.600 237.400 135.800 237.600 ;
        RECT 164.200 237.600 214.200 238.000 ;
        RECT 164.200 237.400 214.400 237.600 ;
        RECT 85.600 237.000 135.600 237.400 ;
        RECT 85.400 236.800 135.600 237.000 ;
        RECT 164.400 237.000 214.400 237.400 ;
        RECT 164.400 236.800 214.600 237.000 ;
        RECT 85.400 236.400 135.400 236.800 ;
        RECT 85.200 236.200 135.400 236.400 ;
        RECT 164.600 236.400 214.600 236.800 ;
        RECT 164.600 236.200 214.800 236.400 ;
        RECT 85.200 235.800 135.200 236.200 ;
        RECT 84.900 235.600 135.200 235.800 ;
        RECT 164.800 235.800 214.800 236.200 ;
        RECT 164.800 235.600 215.000 235.800 ;
        RECT 84.900 235.200 135.000 235.600 ;
        RECT 84.700 235.000 135.000 235.200 ;
        RECT 165.000 235.200 215.000 235.600 ;
        RECT 165.000 235.000 215.300 235.200 ;
        RECT 84.700 234.600 134.700 235.000 ;
        RECT 84.500 234.400 134.700 234.600 ;
        RECT 165.300 234.600 215.300 235.000 ;
        RECT 165.300 234.400 215.500 234.600 ;
        RECT 84.500 234.000 134.500 234.400 ;
        RECT 84.300 233.800 134.500 234.000 ;
        RECT 165.500 234.000 215.500 234.400 ;
        RECT 165.500 233.800 215.700 234.000 ;
        RECT 84.300 233.400 134.300 233.800 ;
        RECT 84.000 233.200 134.300 233.400 ;
        RECT 165.700 233.400 215.700 233.800 ;
        RECT 165.700 233.200 216.000 233.400 ;
        RECT 84.000 232.800 134.000 233.200 ;
        RECT 83.800 232.600 134.000 232.800 ;
        RECT 166.000 232.800 216.000 233.200 ;
        RECT 166.000 232.600 216.200 232.800 ;
        RECT 83.800 232.200 133.800 232.600 ;
        RECT 83.600 232.000 133.800 232.200 ;
        RECT 166.200 232.200 216.200 232.600 ;
        RECT 166.200 232.000 216.400 232.200 ;
        RECT 83.600 231.600 133.600 232.000 ;
        RECT 83.400 231.400 133.600 231.600 ;
        RECT 166.400 231.600 216.400 232.000 ;
        RECT 166.400 231.400 216.600 231.600 ;
        RECT 83.400 231.000 133.400 231.400 ;
        RECT 83.200 230.800 133.400 231.000 ;
        RECT 166.600 231.000 216.600 231.400 ;
        RECT 166.600 230.800 216.800 231.000 ;
        RECT 83.200 230.400 133.200 230.800 ;
        RECT 82.900 230.200 133.200 230.400 ;
        RECT 166.800 230.400 216.800 230.800 ;
        RECT 166.800 230.200 217.100 230.400 ;
        RECT 82.900 229.800 132.900 230.200 ;
        RECT 82.700 229.600 132.900 229.800 ;
        RECT 167.100 229.800 217.100 230.200 ;
        RECT 167.100 229.600 217.300 229.800 ;
        RECT 82.700 229.200 132.700 229.600 ;
        RECT 82.500 229.000 132.700 229.200 ;
        RECT 167.300 229.200 217.300 229.600 ;
        RECT 167.300 229.000 217.500 229.200 ;
        RECT 82.500 228.600 132.500 229.000 ;
        RECT 82.200 228.400 132.500 228.600 ;
        RECT 167.500 228.600 217.500 229.000 ;
        RECT 167.500 228.400 217.800 228.600 ;
        RECT 82.200 228.000 132.200 228.400 ;
        RECT 82.000 227.800 132.200 228.000 ;
        RECT 167.800 228.000 217.800 228.400 ;
        RECT 167.800 227.800 218.000 228.000 ;
        RECT 82.000 227.400 132.000 227.800 ;
        RECT 81.800 227.200 132.000 227.400 ;
        RECT 168.000 227.400 218.000 227.800 ;
        RECT 168.000 227.200 218.200 227.400 ;
        RECT 81.800 226.800 131.800 227.200 ;
        RECT 81.600 226.600 131.800 226.800 ;
        RECT 168.200 226.800 218.200 227.200 ;
        RECT 168.200 226.600 218.400 226.800 ;
        RECT 81.600 226.200 131.600 226.600 ;
        RECT 81.400 226.000 131.600 226.200 ;
        RECT 168.400 226.200 218.400 226.600 ;
        RECT 168.400 226.000 218.600 226.200 ;
        RECT 81.400 225.600 131.400 226.000 ;
        RECT 81.100 225.400 131.400 225.600 ;
        RECT 168.600 225.600 218.600 226.000 ;
        RECT 168.600 225.400 218.900 225.600 ;
        RECT 81.100 225.000 131.100 225.400 ;
        RECT 80.900 224.800 131.100 225.000 ;
        RECT 168.900 225.000 218.900 225.400 ;
        RECT 168.900 224.800 219.100 225.000 ;
        RECT 80.900 224.400 130.900 224.800 ;
        RECT 80.700 224.200 130.900 224.400 ;
        RECT 169.100 224.400 219.100 224.800 ;
        RECT 169.100 224.200 219.300 224.400 ;
        RECT 80.700 223.800 130.700 224.200 ;
        RECT 80.400 223.600 130.700 223.800 ;
        RECT 169.300 223.800 219.300 224.200 ;
        RECT 169.300 223.600 219.600 223.800 ;
        RECT 80.400 223.200 130.400 223.600 ;
        RECT 80.200 223.000 130.400 223.200 ;
        RECT 169.600 223.200 219.600 223.600 ;
        RECT 169.600 223.000 219.800 223.200 ;
        RECT 80.200 222.600 130.200 223.000 ;
        RECT 80.000 222.400 130.200 222.600 ;
        RECT 169.800 222.600 219.800 223.000 ;
        RECT 169.800 222.400 220.000 222.600 ;
        RECT 80.000 222.000 130.000 222.400 ;
        RECT 79.800 221.800 130.000 222.000 ;
        RECT 170.000 222.000 220.000 222.400 ;
        RECT 170.000 221.800 220.200 222.000 ;
        RECT 79.800 221.400 129.800 221.800 ;
        RECT 79.600 221.200 129.800 221.400 ;
        RECT 170.200 221.400 220.200 221.800 ;
        RECT 170.200 221.200 220.400 221.400 ;
        RECT 79.600 220.800 129.600 221.200 ;
        RECT 79.300 220.600 129.600 220.800 ;
        RECT 170.400 220.800 220.400 221.200 ;
        RECT 170.400 220.600 220.700 220.800 ;
        RECT 79.300 220.200 129.300 220.600 ;
        RECT 79.100 220.000 129.300 220.200 ;
        RECT 170.700 220.200 220.700 220.600 ;
        RECT 170.700 220.000 220.900 220.200 ;
        RECT 79.100 219.600 129.100 220.000 ;
        RECT 78.900 219.400 129.100 219.600 ;
        RECT 170.900 219.600 220.900 220.000 ;
        RECT 170.900 219.400 221.100 219.600 ;
        RECT 78.900 219.000 128.900 219.400 ;
        RECT 78.600 218.800 128.900 219.000 ;
        RECT 171.100 219.000 221.100 219.400 ;
        RECT 171.100 218.800 221.400 219.000 ;
        RECT 78.600 218.400 128.600 218.800 ;
        RECT 78.400 218.200 128.600 218.400 ;
        RECT 171.400 218.400 221.400 218.800 ;
        RECT 171.400 218.200 221.600 218.400 ;
        RECT 78.400 217.800 128.400 218.200 ;
        RECT 78.200 217.600 128.400 217.800 ;
        RECT 171.600 217.800 221.600 218.200 ;
        RECT 171.600 217.600 221.800 217.800 ;
        RECT 78.200 217.200 128.200 217.600 ;
        RECT 78.000 217.000 128.200 217.200 ;
        RECT 171.800 217.200 221.800 217.600 ;
        RECT 171.800 217.000 222.000 217.200 ;
        RECT 78.000 216.600 128.000 217.000 ;
        RECT 77.800 216.400 128.000 216.600 ;
        RECT 172.000 216.600 222.000 217.000 ;
        RECT 172.000 216.400 222.200 216.600 ;
        RECT 77.800 216.000 127.800 216.400 ;
        RECT 77.500 215.800 127.800 216.000 ;
        RECT 172.200 216.000 222.200 216.400 ;
        RECT 172.200 215.800 222.500 216.000 ;
        RECT 77.500 215.400 127.500 215.800 ;
        RECT 77.300 215.200 127.500 215.400 ;
        RECT 172.500 215.400 222.500 215.800 ;
        RECT 172.500 215.200 222.700 215.400 ;
        RECT 77.300 214.800 127.300 215.200 ;
        RECT 77.100 214.600 127.300 214.800 ;
        RECT 172.700 214.800 222.700 215.200 ;
        RECT 172.700 214.600 222.900 214.800 ;
        RECT 77.100 214.200 127.100 214.600 ;
        RECT 76.800 214.000 127.100 214.200 ;
        RECT 172.900 214.200 222.900 214.600 ;
        RECT 172.900 214.000 223.200 214.200 ;
        RECT 76.800 213.600 126.800 214.000 ;
        RECT 76.600 213.400 126.800 213.600 ;
        RECT 173.200 213.600 223.200 214.000 ;
        RECT 173.200 213.400 223.400 213.600 ;
        RECT 76.600 213.000 126.600 213.400 ;
        RECT 76.400 212.800 126.600 213.000 ;
        RECT 173.400 213.000 223.400 213.400 ;
        RECT 173.400 212.800 223.600 213.000 ;
        RECT 76.400 212.400 126.400 212.800 ;
        RECT 76.200 212.200 126.400 212.400 ;
        RECT 173.600 212.400 223.600 212.800 ;
        RECT 173.600 212.200 223.800 212.400 ;
        RECT 76.200 211.800 126.200 212.200 ;
        RECT 75.900 211.600 126.200 211.800 ;
        RECT 173.800 211.800 223.800 212.200 ;
        RECT 173.800 211.600 224.000 211.800 ;
        RECT 75.900 211.200 125.900 211.600 ;
        RECT 75.700 211.000 125.900 211.200 ;
        RECT 174.000 211.200 224.000 211.600 ;
        RECT 174.000 211.000 224.300 211.200 ;
        RECT 75.700 210.600 125.700 211.000 ;
        RECT 75.500 210.400 125.700 210.600 ;
        RECT 174.300 210.600 224.300 211.000 ;
        RECT 174.300 210.400 224.500 210.600 ;
        RECT 75.500 210.000 125.500 210.400 ;
        RECT 75.300 209.800 125.500 210.000 ;
        RECT 174.500 210.000 224.500 210.400 ;
        RECT 174.500 209.800 224.700 210.000 ;
        RECT 75.300 209.400 125.300 209.800 ;
        RECT 75.000 209.200 125.300 209.400 ;
        RECT 174.700 209.400 224.700 209.800 ;
        RECT 174.700 209.200 225.000 209.400 ;
        RECT 75.000 208.800 125.000 209.200 ;
        RECT 74.800 208.600 125.000 208.800 ;
        RECT 175.000 208.800 225.000 209.200 ;
        RECT 175.000 208.600 225.200 208.800 ;
        RECT 74.800 208.200 124.800 208.600 ;
        RECT 74.600 208.000 124.800 208.200 ;
        RECT 175.200 208.200 225.200 208.600 ;
        RECT 175.200 208.000 225.400 208.200 ;
        RECT 74.600 207.600 124.600 208.000 ;
        RECT 74.400 207.400 124.600 207.600 ;
        RECT 175.400 207.600 225.400 208.000 ;
        RECT 175.400 207.400 225.600 207.600 ;
        RECT 74.400 207.000 124.400 207.400 ;
        RECT 74.200 206.800 124.400 207.000 ;
        RECT 175.600 207.000 225.600 207.400 ;
        RECT 175.600 206.800 225.800 207.000 ;
        RECT 74.200 206.400 124.200 206.800 ;
        RECT 73.900 206.200 124.200 206.400 ;
        RECT 175.800 206.400 225.800 206.800 ;
        RECT 175.800 206.200 226.100 206.400 ;
        RECT 73.900 205.800 123.900 206.200 ;
        RECT 73.700 205.600 123.900 205.800 ;
        RECT 176.100 205.800 226.100 206.200 ;
        RECT 176.100 205.600 226.300 205.800 ;
        RECT 73.700 205.200 123.700 205.600 ;
        RECT 73.500 205.000 123.700 205.200 ;
        RECT 176.300 205.200 226.300 205.600 ;
        RECT 176.300 205.000 226.500 205.200 ;
        RECT 73.500 204.600 123.500 205.000 ;
        RECT 73.200 204.400 123.500 204.600 ;
        RECT 176.500 204.600 226.500 205.000 ;
        RECT 176.500 204.400 226.800 204.600 ;
        RECT 73.200 204.000 123.200 204.400 ;
        RECT 73.000 203.800 123.200 204.000 ;
        RECT 176.800 204.000 226.800 204.400 ;
        RECT 176.800 203.800 227.000 204.000 ;
        RECT 73.000 203.400 123.000 203.800 ;
        RECT 72.800 203.200 123.000 203.400 ;
        RECT 177.000 203.400 227.000 203.800 ;
        RECT 177.000 203.200 227.200 203.400 ;
        RECT 72.800 202.800 122.800 203.200 ;
        RECT 72.600 202.600 122.800 202.800 ;
        RECT 177.200 202.800 227.200 203.200 ;
        RECT 177.200 202.600 227.400 202.800 ;
        RECT 72.600 202.200 122.600 202.600 ;
        RECT 72.400 202.000 122.600 202.200 ;
        RECT 177.400 202.200 227.400 202.600 ;
        RECT 177.400 202.000 227.600 202.200 ;
        RECT 72.400 201.600 122.400 202.000 ;
        RECT 72.100 201.400 122.400 201.600 ;
        RECT 177.600 201.600 227.600 202.000 ;
        RECT 177.600 201.400 227.900 201.600 ;
        RECT 72.100 201.000 122.100 201.400 ;
        RECT 71.900 200.800 122.100 201.000 ;
        RECT 177.900 201.000 227.900 201.400 ;
        RECT 177.900 200.800 228.100 201.000 ;
        RECT 71.900 200.400 121.900 200.800 ;
        RECT 71.700 200.200 121.900 200.400 ;
        RECT 178.100 200.400 228.100 200.800 ;
        RECT 178.100 200.200 228.300 200.400 ;
        RECT 71.700 199.800 121.700 200.200 ;
        RECT 71.400 199.600 121.700 199.800 ;
        RECT 178.300 199.800 228.300 200.200 ;
        RECT 178.300 199.600 228.600 199.800 ;
        RECT 71.400 199.200 121.400 199.600 ;
        RECT 71.200 199.000 121.400 199.200 ;
        RECT 178.600 199.200 228.600 199.600 ;
        RECT 178.600 199.000 228.800 199.200 ;
        RECT 71.200 198.600 121.200 199.000 ;
        RECT 71.000 198.400 121.200 198.600 ;
        RECT 178.800 198.600 228.800 199.000 ;
        RECT 178.800 198.400 229.000 198.600 ;
        RECT 71.000 198.000 121.000 198.400 ;
        RECT 70.800 197.800 121.000 198.000 ;
        RECT 179.000 198.000 229.000 198.400 ;
        RECT 179.000 197.800 229.200 198.000 ;
        RECT 70.800 197.400 120.800 197.800 ;
        RECT 70.600 197.200 120.800 197.400 ;
        RECT 179.200 197.400 229.200 197.800 ;
        RECT 179.200 197.200 229.400 197.400 ;
        RECT 70.600 196.800 120.600 197.200 ;
        RECT 70.300 196.600 120.600 196.800 ;
        RECT 179.400 196.800 229.400 197.200 ;
        RECT 179.400 196.600 229.700 196.800 ;
        RECT 70.300 196.200 120.300 196.600 ;
        RECT 70.100 196.000 120.300 196.200 ;
        RECT 179.700 196.200 229.700 196.600 ;
        RECT 179.700 196.000 229.900 196.200 ;
        RECT 70.100 195.600 120.100 196.000 ;
        RECT 69.900 195.400 120.100 195.600 ;
        RECT 179.900 195.600 229.900 196.000 ;
        RECT 179.900 195.400 230.100 195.600 ;
        RECT 69.900 195.000 119.900 195.400 ;
        RECT 69.600 194.800 119.900 195.000 ;
        RECT 180.100 195.000 230.100 195.400 ;
        RECT 180.100 194.800 230.400 195.000 ;
        RECT 69.600 194.400 119.600 194.800 ;
        RECT 69.400 194.200 119.600 194.400 ;
        RECT 180.400 194.400 230.400 194.800 ;
        RECT 180.400 194.200 230.600 194.400 ;
        RECT 69.400 193.800 119.400 194.200 ;
        RECT 69.200 193.600 119.400 193.800 ;
        RECT 180.600 193.800 230.600 194.200 ;
        RECT 180.600 193.600 230.800 193.800 ;
        RECT 69.200 193.200 119.200 193.600 ;
        RECT 69.000 193.000 119.200 193.200 ;
        RECT 180.800 193.200 230.800 193.600 ;
        RECT 180.800 193.000 231.000 193.200 ;
        RECT 69.000 192.600 119.000 193.000 ;
        RECT 68.800 192.400 119.000 192.600 ;
        RECT 181.000 192.600 231.000 193.000 ;
        RECT 181.000 192.400 231.200 192.600 ;
        RECT 68.800 192.000 118.800 192.400 ;
        RECT 68.500 191.800 118.800 192.000 ;
        RECT 181.200 192.000 231.200 192.400 ;
        RECT 181.200 191.800 231.500 192.000 ;
        RECT 68.500 191.400 118.500 191.800 ;
        RECT 68.300 191.200 118.500 191.400 ;
        RECT 181.500 191.400 231.500 191.800 ;
        RECT 181.500 191.200 231.700 191.400 ;
        RECT 68.300 190.800 118.300 191.200 ;
        RECT 68.100 190.600 118.300 190.800 ;
        RECT 181.700 190.800 231.700 191.200 ;
        RECT 181.700 190.600 231.900 190.800 ;
        RECT 68.100 190.200 118.100 190.600 ;
        RECT 67.800 190.000 118.100 190.200 ;
        RECT 181.900 190.200 231.900 190.600 ;
        RECT 181.900 190.000 232.200 190.200 ;
        RECT 67.800 189.600 117.800 190.000 ;
        RECT 67.600 189.400 117.800 189.600 ;
        RECT 182.200 189.600 232.200 190.000 ;
        RECT 182.200 189.400 232.400 189.600 ;
        RECT 67.600 189.000 117.600 189.400 ;
        RECT 67.400 188.800 117.600 189.000 ;
        RECT 182.400 189.000 232.400 189.400 ;
        RECT 182.400 188.800 232.600 189.000 ;
        RECT 67.400 188.400 117.400 188.800 ;
        RECT 67.200 188.200 117.400 188.400 ;
        RECT 182.600 188.400 232.600 188.800 ;
        RECT 182.600 188.200 232.800 188.400 ;
        RECT 67.200 187.800 117.200 188.200 ;
        RECT 66.900 187.600 117.200 187.800 ;
        RECT 182.800 187.800 232.800 188.200 ;
        RECT 182.800 187.600 233.000 187.800 ;
        RECT 66.900 187.200 116.900 187.600 ;
        RECT 66.700 187.000 116.900 187.200 ;
        RECT 183.000 187.200 233.000 187.600 ;
        RECT 183.000 187.000 233.300 187.200 ;
        RECT 66.700 186.600 116.700 187.000 ;
        RECT 66.500 186.400 116.700 186.600 ;
        RECT 183.300 186.600 233.300 187.000 ;
        RECT 183.300 186.400 233.500 186.600 ;
        RECT 66.500 186.000 116.500 186.400 ;
        RECT 66.300 185.800 116.500 186.000 ;
        RECT 183.500 186.000 233.500 186.400 ;
        RECT 183.500 185.800 233.700 186.000 ;
        RECT 66.300 185.400 116.300 185.800 ;
        RECT 66.000 185.200 116.300 185.400 ;
        RECT 183.700 185.400 233.700 185.800 ;
        RECT 183.700 185.200 234.000 185.400 ;
        RECT 66.000 184.800 116.000 185.200 ;
        RECT 65.800 184.600 116.000 184.800 ;
        RECT 184.000 184.800 234.000 185.200 ;
        RECT 184.000 184.600 234.200 184.800 ;
        RECT 65.800 184.200 115.800 184.600 ;
        RECT 65.600 184.000 115.800 184.200 ;
        RECT 184.200 184.200 234.200 184.600 ;
        RECT 184.200 184.000 234.400 184.200 ;
        RECT 65.600 183.600 115.600 184.000 ;
        RECT 65.400 183.400 115.600 183.600 ;
        RECT 184.400 183.600 234.400 184.000 ;
        RECT 184.400 183.400 234.600 183.600 ;
        RECT 65.400 183.000 115.400 183.400 ;
        RECT 65.200 182.800 115.400 183.000 ;
        RECT 184.600 183.000 234.600 183.400 ;
        RECT 184.600 182.800 234.800 183.000 ;
        RECT 65.200 182.400 115.200 182.800 ;
        RECT 64.900 182.200 115.200 182.400 ;
        RECT 184.800 182.400 234.800 182.800 ;
        RECT 184.800 182.200 235.100 182.400 ;
        RECT 64.900 181.800 114.900 182.200 ;
        RECT 64.700 181.600 114.900 181.800 ;
        RECT 185.100 181.800 235.100 182.200 ;
        RECT 185.100 181.600 235.300 181.800 ;
        RECT 64.700 181.200 114.700 181.600 ;
        RECT 64.500 181.000 114.700 181.200 ;
        RECT 185.300 181.200 235.300 181.600 ;
        RECT 185.300 181.000 235.500 181.200 ;
        RECT 64.500 180.600 114.500 181.000 ;
        RECT 64.200 180.400 114.500 180.600 ;
        RECT 185.500 180.600 235.500 181.000 ;
        RECT 185.500 180.400 235.800 180.600 ;
        RECT 64.200 180.000 114.200 180.400 ;
        RECT 64.000 179.800 114.200 180.000 ;
        RECT 185.800 180.000 235.800 180.400 ;
        RECT 185.800 179.800 236.000 180.000 ;
        RECT 64.000 179.400 114.000 179.800 ;
        RECT 63.800 179.200 114.000 179.400 ;
        RECT 186.000 179.400 236.000 179.800 ;
        RECT 186.000 179.200 236.200 179.400 ;
        RECT 63.800 178.800 113.800 179.200 ;
        RECT 63.600 178.600 113.800 178.800 ;
        RECT 186.200 178.800 236.200 179.200 ;
        RECT 186.200 178.600 236.400 178.800 ;
        RECT 63.600 178.200 113.600 178.600 ;
        RECT 63.300 178.000 113.600 178.200 ;
        RECT 186.400 178.200 236.400 178.600 ;
        RECT 186.400 178.000 236.600 178.200 ;
        RECT 63.300 177.600 113.400 178.000 ;
        RECT 63.100 177.400 113.400 177.600 ;
        RECT 186.600 177.600 236.600 178.000 ;
        RECT 186.600 177.400 236.900 177.600 ;
        RECT 63.100 177.000 113.100 177.400 ;
        RECT 62.900 176.800 113.100 177.000 ;
        RECT 186.900 177.000 236.900 177.400 ;
        RECT 186.900 176.800 237.100 177.000 ;
        RECT 62.900 176.400 112.900 176.800 ;
        RECT 62.700 176.200 112.900 176.400 ;
        RECT 187.100 176.400 237.100 176.800 ;
        RECT 187.100 176.200 237.300 176.400 ;
        RECT 62.700 175.800 112.700 176.200 ;
        RECT 62.400 175.600 112.700 175.800 ;
        RECT 187.300 175.800 237.300 176.200 ;
        RECT 187.300 175.600 237.600 175.800 ;
        RECT 62.400 175.200 112.400 175.600 ;
        RECT 62.200 175.000 112.400 175.200 ;
        RECT 187.600 175.200 237.600 175.600 ;
        RECT 187.600 175.000 237.800 175.200 ;
        RECT 62.200 174.600 112.200 175.000 ;
        RECT 62.000 174.400 112.200 174.600 ;
        RECT 187.800 174.600 237.800 175.000 ;
        RECT 187.800 174.400 238.000 174.600 ;
        RECT 62.000 174.000 112.000 174.400 ;
        RECT 61.800 173.800 112.000 174.000 ;
        RECT 188.000 174.000 238.000 174.400 ;
        RECT 188.000 173.800 238.200 174.000 ;
        RECT 61.800 173.400 111.800 173.800 ;
        RECT 61.600 173.200 111.800 173.400 ;
        RECT 188.200 173.400 238.200 173.800 ;
        RECT 188.200 173.200 238.400 173.400 ;
        RECT 61.600 172.800 111.600 173.200 ;
        RECT 61.300 172.600 111.600 172.800 ;
        RECT 188.400 172.800 238.400 173.200 ;
        RECT 188.400 172.600 238.700 172.800 ;
        RECT 61.300 172.200 111.300 172.600 ;
        RECT 61.100 172.000 111.300 172.200 ;
        RECT 188.700 172.200 238.700 172.600 ;
        RECT 188.700 172.000 238.900 172.200 ;
        RECT 61.100 171.600 111.100 172.000 ;
        RECT 60.900 171.400 111.100 171.600 ;
        RECT 188.900 171.600 238.900 172.000 ;
        RECT 188.900 171.400 239.100 171.600 ;
        RECT 60.900 171.000 110.900 171.400 ;
        RECT 60.600 170.800 110.900 171.000 ;
        RECT 189.100 171.000 239.100 171.400 ;
        RECT 189.100 170.800 239.400 171.000 ;
        RECT 60.600 170.400 110.600 170.800 ;
        RECT 60.400 170.200 110.600 170.400 ;
        RECT 189.400 170.400 239.400 170.800 ;
        RECT 189.400 170.200 239.600 170.400 ;
        RECT 60.400 169.800 110.400 170.200 ;
        RECT 60.200 169.600 110.400 169.800 ;
        RECT 189.600 169.800 239.600 170.200 ;
        RECT 189.600 169.600 239.800 169.800 ;
        RECT 60.200 169.200 110.200 169.600 ;
        RECT 60.000 169.000 110.200 169.200 ;
        RECT 189.800 169.200 239.800 169.600 ;
        RECT 189.800 169.000 240.000 169.200 ;
        RECT 60.000 168.600 110.000 169.000 ;
        RECT 59.800 168.400 110.000 168.600 ;
        RECT 190.000 168.600 240.000 169.000 ;
        RECT 190.000 168.400 240.200 168.600 ;
        RECT 59.800 168.000 109.800 168.400 ;
        RECT 59.500 167.800 109.800 168.000 ;
        RECT 190.200 168.000 240.200 168.400 ;
        RECT 190.200 167.800 240.500 168.000 ;
        RECT 59.500 167.400 109.500 167.800 ;
        RECT 59.300 167.200 109.500 167.400 ;
        RECT 190.500 167.400 240.500 167.800 ;
        RECT 190.500 167.200 240.700 167.400 ;
        RECT 59.300 166.800 109.300 167.200 ;
        RECT 59.100 166.600 109.300 166.800 ;
        RECT 190.700 166.800 240.700 167.200 ;
        RECT 190.700 166.600 240.900 166.800 ;
        RECT 59.100 166.200 109.100 166.600 ;
        RECT 58.800 166.000 109.100 166.200 ;
        RECT 190.900 166.200 240.900 166.600 ;
        RECT 190.900 166.000 241.200 166.200 ;
        RECT 58.800 165.600 108.800 166.000 ;
        RECT 58.600 165.400 108.800 165.600 ;
        RECT 191.200 165.600 241.200 166.000 ;
        RECT 191.200 165.400 241.400 165.600 ;
        RECT 58.600 165.000 108.600 165.400 ;
        RECT 58.400 164.800 108.600 165.000 ;
        RECT 191.400 165.000 241.400 165.400 ;
        RECT 191.400 164.800 241.600 165.000 ;
        RECT 58.400 164.400 108.400 164.800 ;
        RECT 58.200 164.200 108.400 164.400 ;
        RECT 191.600 164.400 241.600 164.800 ;
        RECT 191.600 164.200 241.800 164.400 ;
        RECT 58.200 163.800 108.200 164.200 ;
        RECT 58.000 163.600 108.200 163.800 ;
        RECT 191.800 163.800 241.800 164.200 ;
        RECT 191.800 163.600 242.000 163.800 ;
        RECT 58.000 163.200 108.000 163.600 ;
        RECT 57.700 163.000 108.000 163.200 ;
        RECT 192.000 163.200 242.000 163.600 ;
        RECT 192.000 163.000 242.300 163.200 ;
        RECT 57.700 162.600 107.700 163.000 ;
        RECT 57.500 162.400 107.700 162.600 ;
        RECT 192.300 162.600 242.300 163.000 ;
        RECT 192.300 162.400 242.500 162.600 ;
        RECT 57.500 162.000 107.500 162.400 ;
        RECT 192.500 162.000 242.500 162.400 ;
        RECT 57.300 161.400 242.700 162.000 ;
        RECT 57.000 160.800 243.000 161.400 ;
        RECT 56.800 160.200 243.200 160.800 ;
        RECT 56.600 159.600 243.400 160.200 ;
        RECT 56.400 159.000 243.600 159.600 ;
        RECT 56.100 158.400 243.900 159.000 ;
        RECT 55.900 157.800 244.100 158.400 ;
        RECT 55.700 157.200 244.300 157.800 ;
        RECT 55.500 156.600 244.500 157.200 ;
        RECT 55.200 156.000 244.800 156.600 ;
        RECT 55.000 155.400 245.000 156.000 ;
        RECT 54.800 154.800 245.200 155.400 ;
        RECT 54.600 154.200 245.400 154.800 ;
        RECT 54.300 153.600 245.600 154.200 ;
        RECT 54.100 153.000 245.900 153.600 ;
        RECT 53.900 152.400 246.100 153.000 ;
        RECT 53.700 151.800 246.300 152.400 ;
        RECT 53.400 151.200 246.600 151.800 ;
        RECT 53.200 150.600 246.800 151.200 ;
        RECT 53.000 150.000 247.000 150.600 ;
        RECT 52.800 149.400 247.200 150.000 ;
        RECT 52.600 148.800 247.400 149.400 ;
        RECT 52.300 148.200 247.700 148.800 ;
        RECT 52.100 147.600 247.900 148.200 ;
        RECT 51.900 147.000 248.100 147.600 ;
        RECT 51.600 146.400 248.400 147.000 ;
        RECT 51.400 145.800 248.600 146.400 ;
        RECT 51.200 145.200 248.800 145.800 ;
        RECT 51.000 144.600 249.000 145.200 ;
        RECT 50.800 144.000 249.200 144.600 ;
        RECT 50.500 143.400 249.500 144.000 ;
        RECT 50.300 142.800 249.700 143.400 ;
        RECT 50.100 142.200 249.900 142.800 ;
        RECT 49.800 141.600 250.200 142.200 ;
        RECT 49.600 141.000 250.400 141.600 ;
        RECT 49.400 140.400 250.600 141.000 ;
        RECT 49.200 139.800 250.800 140.400 ;
        RECT 49.000 139.200 251.000 139.800 ;
        RECT 48.700 138.600 251.300 139.200 ;
        RECT 48.500 138.000 251.500 138.600 ;
        RECT 48.300 137.400 251.700 138.000 ;
        RECT 48.000 136.800 252.000 137.400 ;
        RECT 47.800 136.200 252.200 136.800 ;
        RECT 47.600 135.600 252.400 136.200 ;
        RECT 47.400 135.000 252.600 135.600 ;
        RECT 47.100 134.400 252.900 135.000 ;
        RECT 46.900 133.800 253.100 134.400 ;
        RECT 46.700 133.200 253.300 133.800 ;
        RECT 46.500 132.600 253.500 133.200 ;
        RECT 46.200 132.000 253.800 132.600 ;
        RECT 46.000 131.400 254.000 132.000 ;
        RECT 45.800 130.800 254.200 131.400 ;
        RECT 45.600 130.200 254.400 130.800 ;
        RECT 45.300 129.600 254.600 130.200 ;
        RECT 45.100 129.000 254.900 129.600 ;
        RECT 44.900 128.400 255.100 129.000 ;
        RECT 44.700 127.800 255.300 128.400 ;
        RECT 44.400 127.200 255.600 127.800 ;
        RECT 44.200 126.600 255.800 127.200 ;
        RECT 44.000 126.000 256.000 126.600 ;
        RECT 43.800 125.400 256.200 126.000 ;
        RECT 43.600 124.800 256.400 125.400 ;
        RECT 43.300 124.200 256.700 124.800 ;
        RECT 43.100 123.600 256.900 124.200 ;
        RECT 42.900 123.000 257.100 123.600 ;
        RECT 42.600 122.400 257.400 123.000 ;
        RECT 42.400 122.200 257.600 122.400 ;
        RECT 42.400 121.800 92.400 122.200 ;
        RECT 42.200 121.600 92.400 121.800 ;
        RECT 207.600 121.800 257.600 122.200 ;
        RECT 207.600 121.600 257.800 121.800 ;
        RECT 42.200 121.200 92.200 121.600 ;
        RECT 42.000 121.000 92.200 121.200 ;
        RECT 207.800 121.200 257.800 121.600 ;
        RECT 207.800 121.000 258.000 121.200 ;
        RECT 42.000 120.600 92.000 121.000 ;
        RECT 41.800 120.400 92.000 120.600 ;
        RECT 208.000 120.600 258.000 121.000 ;
        RECT 208.000 120.400 258.200 120.600 ;
        RECT 41.800 120.000 91.800 120.400 ;
        RECT 41.500 119.800 91.800 120.000 ;
        RECT 208.200 120.000 258.200 120.400 ;
        RECT 208.200 119.800 258.500 120.000 ;
        RECT 41.500 119.400 91.500 119.800 ;
        RECT 41.300 119.200 91.500 119.400 ;
        RECT 208.500 119.400 258.500 119.800 ;
        RECT 208.500 119.200 258.700 119.400 ;
        RECT 41.300 118.800 91.300 119.200 ;
        RECT 41.100 118.600 91.300 118.800 ;
        RECT 208.700 118.800 258.700 119.200 ;
        RECT 208.700 118.600 258.900 118.800 ;
        RECT 41.100 118.200 91.100 118.600 ;
        RECT 40.800 118.000 91.100 118.200 ;
        RECT 208.900 118.200 258.900 118.600 ;
        RECT 208.900 118.000 259.100 118.200 ;
        RECT 40.800 117.600 90.800 118.000 ;
        RECT 40.600 117.400 90.800 117.600 ;
        RECT 209.200 117.600 259.100 118.000 ;
        RECT 209.200 117.400 259.400 117.600 ;
        RECT 40.600 117.000 90.600 117.400 ;
        RECT 40.400 116.800 90.600 117.000 ;
        RECT 209.400 117.000 259.400 117.400 ;
        RECT 209.400 116.800 259.600 117.000 ;
        RECT 40.400 116.400 90.400 116.800 ;
        RECT 40.200 116.200 90.400 116.400 ;
        RECT 209.600 116.400 259.600 116.800 ;
        RECT 209.600 116.200 259.800 116.400 ;
        RECT 40.200 115.800 90.200 116.200 ;
        RECT 40.000 115.600 90.200 115.800 ;
        RECT 209.800 115.800 259.800 116.200 ;
        RECT 209.800 115.600 260.000 115.800 ;
        RECT 40.000 115.200 90.000 115.600 ;
        RECT 39.700 115.000 90.000 115.200 ;
        RECT 210.000 115.200 260.000 115.600 ;
        RECT 210.000 115.000 260.300 115.200 ;
        RECT 39.700 114.600 89.700 115.000 ;
        RECT 39.500 114.400 89.700 114.600 ;
        RECT 210.300 114.600 260.300 115.000 ;
        RECT 210.300 114.400 260.500 114.600 ;
        RECT 39.500 114.000 89.500 114.400 ;
        RECT 39.300 113.800 89.500 114.000 ;
        RECT 210.500 114.000 260.500 114.400 ;
        RECT 210.500 113.800 260.700 114.000 ;
        RECT 39.300 113.400 89.300 113.800 ;
        RECT 39.000 113.200 89.300 113.400 ;
        RECT 210.700 113.400 260.700 113.800 ;
        RECT 210.700 113.200 261.000 113.400 ;
        RECT 39.000 112.800 89.000 113.200 ;
        RECT 38.800 112.600 89.000 112.800 ;
        RECT 211.000 112.800 261.000 113.200 ;
        RECT 211.000 112.600 261.200 112.800 ;
        RECT 38.800 112.200 88.800 112.600 ;
        RECT 38.600 112.000 88.800 112.200 ;
        RECT 211.200 112.200 261.200 112.600 ;
        RECT 211.200 112.000 261.400 112.200 ;
        RECT 38.600 111.600 88.600 112.000 ;
        RECT 38.400 111.400 88.600 111.600 ;
        RECT 211.400 111.600 261.400 112.000 ;
        RECT 211.400 111.400 261.600 111.600 ;
        RECT 38.400 111.000 88.400 111.400 ;
        RECT 38.100 110.800 88.400 111.000 ;
        RECT 211.600 111.000 261.600 111.400 ;
        RECT 211.600 110.800 261.900 111.000 ;
        RECT 38.100 110.400 88.100 110.800 ;
        RECT 37.900 110.200 88.100 110.400 ;
        RECT 211.900 110.400 261.900 110.800 ;
        RECT 211.900 110.200 262.100 110.400 ;
        RECT 37.900 109.800 87.900 110.200 ;
        RECT 37.700 109.600 87.900 109.800 ;
        RECT 212.100 109.800 262.100 110.200 ;
        RECT 212.100 109.600 262.300 109.800 ;
        RECT 37.700 109.200 87.700 109.600 ;
        RECT 37.500 109.000 87.700 109.200 ;
        RECT 212.300 109.200 262.300 109.600 ;
        RECT 212.300 109.000 262.500 109.200 ;
        RECT 37.500 108.600 87.500 109.000 ;
        RECT 37.200 108.400 87.500 108.600 ;
        RECT 212.500 108.600 262.500 109.000 ;
        RECT 212.500 108.400 262.800 108.600 ;
        RECT 37.200 108.000 87.200 108.400 ;
        RECT 37.000 107.800 87.200 108.000 ;
        RECT 212.800 108.000 262.800 108.400 ;
        RECT 212.800 107.800 263.000 108.000 ;
        RECT 37.000 107.400 87.000 107.800 ;
        RECT 36.800 107.200 87.000 107.400 ;
        RECT 213.000 107.400 263.000 107.800 ;
        RECT 213.000 107.200 263.200 107.400 ;
        RECT 36.800 106.800 86.800 107.200 ;
        RECT 36.600 106.600 86.800 106.800 ;
        RECT 213.200 106.800 263.200 107.200 ;
        RECT 213.200 106.600 263.400 106.800 ;
        RECT 36.600 106.200 86.600 106.600 ;
        RECT 36.300 106.000 86.600 106.200 ;
        RECT 213.400 106.200 263.400 106.600 ;
        RECT 213.400 106.000 263.600 106.200 ;
        RECT 36.300 105.600 86.400 106.000 ;
        RECT 36.100 105.400 86.400 105.600 ;
        RECT 213.600 105.600 263.600 106.000 ;
        RECT 213.600 105.400 263.900 105.600 ;
        RECT 36.100 105.000 86.100 105.400 ;
        RECT 35.900 104.800 86.100 105.000 ;
        RECT 213.900 105.000 263.900 105.400 ;
        RECT 213.900 104.800 264.100 105.000 ;
        RECT 35.900 104.400 85.900 104.800 ;
        RECT 35.700 104.200 85.900 104.400 ;
        RECT 214.100 104.400 264.100 104.800 ;
        RECT 214.100 104.200 264.300 104.400 ;
        RECT 35.700 103.800 85.700 104.200 ;
        RECT 35.400 103.600 85.700 103.800 ;
        RECT 214.300 103.800 264.300 104.200 ;
        RECT 214.300 103.600 264.600 103.800 ;
        RECT 35.400 103.200 85.400 103.600 ;
        RECT 35.200 103.000 85.400 103.200 ;
        RECT 214.600 103.200 264.600 103.600 ;
        RECT 214.600 103.000 264.800 103.200 ;
        RECT 35.200 102.600 85.200 103.000 ;
        RECT 35.000 102.400 85.200 102.600 ;
        RECT 214.800 102.600 264.800 103.000 ;
        RECT 214.800 102.400 265.000 102.600 ;
        RECT 35.000 102.000 85.000 102.400 ;
        RECT 34.800 101.800 85.000 102.000 ;
        RECT 215.000 102.000 265.000 102.400 ;
        RECT 215.000 101.800 265.200 102.000 ;
        RECT 34.800 101.400 84.800 101.800 ;
        RECT 34.600 101.200 84.800 101.400 ;
        RECT 215.200 101.400 265.200 101.800 ;
        RECT 215.200 101.200 265.400 101.400 ;
        RECT 34.600 100.800 84.600 101.200 ;
        RECT 34.300 100.600 84.600 100.800 ;
        RECT 215.400 100.800 265.400 101.200 ;
        RECT 215.400 100.600 265.700 100.800 ;
        RECT 34.300 100.200 84.300 100.600 ;
        RECT 34.100 100.000 84.300 100.200 ;
        RECT 215.700 100.200 265.700 100.600 ;
        RECT 215.700 100.000 265.900 100.200 ;
        RECT 34.100 99.600 84.100 100.000 ;
        RECT 33.900 99.400 84.100 99.600 ;
        RECT 215.900 99.600 265.900 100.000 ;
        RECT 215.900 99.400 266.100 99.600 ;
        RECT 33.900 99.000 83.900 99.400 ;
        RECT 33.600 98.800 83.900 99.000 ;
        RECT 216.100 99.000 266.100 99.400 ;
        RECT 216.100 98.800 266.400 99.000 ;
        RECT 33.600 98.400 83.600 98.800 ;
        RECT 33.400 98.200 83.600 98.400 ;
        RECT 216.400 98.400 266.400 98.800 ;
        RECT 216.400 98.200 266.600 98.400 ;
        RECT 33.400 97.800 83.400 98.200 ;
        RECT 33.200 97.600 83.400 97.800 ;
        RECT 216.600 97.800 266.600 98.200 ;
        RECT 216.600 97.600 266.800 97.800 ;
        RECT 33.200 97.200 83.200 97.600 ;
        RECT 33.000 97.000 83.200 97.200 ;
        RECT 216.800 97.200 266.800 97.600 ;
        RECT 216.800 97.000 267.000 97.200 ;
        RECT 33.000 96.600 83.000 97.000 ;
        RECT 32.800 96.400 83.000 96.600 ;
        RECT 217.000 96.600 267.000 97.000 ;
        RECT 217.000 96.400 267.200 96.600 ;
        RECT 32.800 96.000 82.800 96.400 ;
        RECT 32.500 95.800 82.800 96.000 ;
        RECT 217.200 96.000 267.200 96.400 ;
        RECT 217.200 95.800 267.500 96.000 ;
        RECT 32.500 95.400 82.500 95.800 ;
        RECT 32.300 95.200 82.500 95.400 ;
        RECT 217.500 95.400 267.500 95.800 ;
        RECT 217.500 95.200 267.700 95.400 ;
        RECT 32.300 94.800 82.300 95.200 ;
        RECT 32.100 94.600 82.300 94.800 ;
        RECT 217.700 94.800 267.700 95.200 ;
        RECT 217.700 94.600 267.900 94.800 ;
        RECT 32.100 94.200 82.100 94.600 ;
        RECT 31.800 94.000 82.100 94.200 ;
        RECT 217.900 94.200 267.900 94.600 ;
        RECT 217.900 94.000 268.200 94.200 ;
        RECT 31.800 93.600 81.800 94.000 ;
        RECT 31.600 93.400 81.800 93.600 ;
        RECT 218.200 93.600 268.200 94.000 ;
        RECT 218.200 93.400 268.400 93.600 ;
        RECT 31.600 93.000 81.600 93.400 ;
        RECT 31.400 92.800 81.600 93.000 ;
        RECT 218.400 93.000 268.400 93.400 ;
        RECT 218.400 92.800 268.600 93.000 ;
        RECT 31.400 92.400 81.400 92.800 ;
        RECT 31.200 92.200 81.400 92.400 ;
        RECT 218.600 92.400 268.600 92.800 ;
        RECT 218.600 92.200 268.800 92.400 ;
        RECT 31.200 91.800 81.200 92.200 ;
        RECT 31.000 91.600 81.200 91.800 ;
        RECT 218.800 91.800 268.800 92.200 ;
        RECT 218.800 91.600 269.000 91.800 ;
        RECT 31.000 91.200 81.000 91.600 ;
        RECT 30.700 91.000 81.000 91.200 ;
        RECT 219.000 91.200 269.000 91.600 ;
        RECT 219.000 91.000 269.300 91.200 ;
        RECT 30.700 90.600 80.700 91.000 ;
        RECT 30.500 90.400 80.700 90.600 ;
        RECT 219.300 90.600 269.300 91.000 ;
        RECT 219.300 90.400 269.500 90.600 ;
        RECT 30.500 90.000 80.500 90.400 ;
        RECT 30.300 89.800 80.500 90.000 ;
        RECT 219.500 90.000 269.500 90.400 ;
        RECT 219.500 89.800 269.700 90.000 ;
        RECT 30.300 89.400 80.300 89.800 ;
        RECT 30.000 89.200 80.300 89.400 ;
        RECT 219.700 89.400 269.700 89.800 ;
        RECT 219.700 89.200 270.000 89.400 ;
        RECT 30.000 88.800 80.000 89.200 ;
        RECT 29.800 88.600 80.000 88.800 ;
        RECT 220.000 88.800 270.000 89.200 ;
        RECT 220.000 88.600 270.200 88.800 ;
        RECT 29.800 88.200 79.800 88.600 ;
        RECT 29.600 88.000 79.800 88.200 ;
        RECT 220.200 88.200 270.200 88.600 ;
        RECT 220.200 88.000 270.400 88.200 ;
        RECT 29.600 87.600 79.600 88.000 ;
        RECT 29.400 87.400 79.600 87.600 ;
        RECT 220.400 87.600 270.400 88.000 ;
        RECT 220.400 87.400 270.600 87.600 ;
        RECT 29.400 87.000 79.400 87.400 ;
        RECT 29.100 86.800 79.400 87.000 ;
        RECT 220.600 87.000 270.600 87.400 ;
        RECT 220.600 86.800 270.800 87.000 ;
        RECT 29.100 86.400 79.100 86.800 ;
        RECT 28.900 86.200 79.100 86.400 ;
        RECT 220.900 86.400 270.800 86.800 ;
        RECT 220.900 86.200 271.100 86.400 ;
        RECT 28.900 85.800 78.900 86.200 ;
        RECT 28.700 85.600 78.900 85.800 ;
        RECT 221.100 85.800 271.100 86.200 ;
        RECT 221.100 85.600 271.300 85.800 ;
        RECT 28.700 85.200 78.700 85.600 ;
        RECT 28.500 85.000 78.700 85.200 ;
        RECT 221.300 85.200 271.300 85.600 ;
        RECT 221.300 85.000 271.500 85.200 ;
        RECT 28.500 84.600 78.500 85.000 ;
        RECT 28.200 84.400 78.500 84.600 ;
        RECT 221.500 84.600 271.500 85.000 ;
        RECT 221.500 84.400 271.800 84.600 ;
        RECT 28.200 84.000 78.200 84.400 ;
        RECT 28.000 83.800 78.200 84.000 ;
        RECT 221.800 84.000 271.800 84.400 ;
        RECT 221.800 83.800 272.000 84.000 ;
        RECT 28.000 83.400 78.000 83.800 ;
        RECT 27.800 83.200 78.000 83.400 ;
        RECT 222.000 83.400 272.000 83.800 ;
        RECT 222.000 83.200 272.200 83.400 ;
        RECT 27.800 82.800 77.800 83.200 ;
        RECT 27.600 82.600 77.800 82.800 ;
        RECT 222.200 82.800 272.200 83.200 ;
        RECT 222.200 82.600 272.400 82.800 ;
        RECT 27.600 82.200 77.600 82.600 ;
        RECT 27.300 82.000 77.600 82.200 ;
        RECT 222.400 82.200 272.400 82.600 ;
        RECT 222.400 82.000 272.600 82.200 ;
        RECT 27.300 81.600 77.400 82.000 ;
        RECT 27.100 81.400 77.400 81.600 ;
        RECT 222.600 81.600 272.600 82.000 ;
        RECT 222.600 81.400 272.900 81.600 ;
        RECT 27.100 81.000 77.100 81.400 ;
        RECT 26.900 80.800 77.100 81.000 ;
        RECT 222.900 81.000 272.900 81.400 ;
        RECT 222.900 80.800 273.100 81.000 ;
        RECT 26.900 80.400 76.900 80.800 ;
        RECT 26.700 80.200 76.900 80.400 ;
        RECT 223.100 80.400 273.100 80.800 ;
        RECT 223.100 80.200 273.300 80.400 ;
        RECT 26.700 79.800 76.700 80.200 ;
        RECT 26.500 79.600 76.700 79.800 ;
        RECT 223.300 79.800 273.300 80.200 ;
        RECT 223.300 79.600 273.600 79.800 ;
        RECT 26.500 79.200 76.400 79.600 ;
        RECT 26.200 79.000 76.400 79.200 ;
        RECT 223.600 79.200 273.600 79.600 ;
        RECT 223.600 79.000 273.800 79.200 ;
        RECT 26.200 78.600 76.200 79.000 ;
        RECT 26.000 78.400 76.200 78.600 ;
        RECT 223.800 78.600 273.800 79.000 ;
        RECT 223.800 78.400 274.000 78.600 ;
        RECT 26.000 78.000 76.000 78.400 ;
        RECT 25.800 77.800 76.000 78.000 ;
        RECT 224.000 78.000 274.000 78.400 ;
        RECT 224.000 77.800 274.200 78.000 ;
        RECT 25.800 77.400 75.800 77.800 ;
        RECT 25.500 77.200 75.800 77.400 ;
        RECT 224.200 77.400 274.200 77.800 ;
        RECT 224.200 77.200 274.400 77.400 ;
        RECT 25.500 76.800 75.600 77.200 ;
        RECT 25.300 76.600 75.600 76.800 ;
        RECT 224.400 76.800 274.400 77.200 ;
        RECT 224.400 76.600 274.700 76.800 ;
        RECT 25.300 76.200 75.300 76.600 ;
        RECT 25.100 76.000 75.300 76.200 ;
        RECT 224.700 76.200 274.700 76.600 ;
        RECT 224.700 76.000 274.900 76.200 ;
        RECT 25.100 75.600 75.100 76.000 ;
        RECT 24.900 75.400 75.100 75.600 ;
        RECT 224.900 75.600 274.900 76.000 ;
        RECT 224.900 75.400 275.100 75.600 ;
        RECT 24.900 75.000 74.900 75.400 ;
        RECT 24.600 74.800 74.900 75.000 ;
        RECT 225.100 75.000 275.100 75.400 ;
        RECT 225.100 74.800 275.400 75.000 ;
        RECT 24.600 74.400 74.600 74.800 ;
        RECT 24.400 74.200 74.600 74.400 ;
        RECT 225.400 74.400 275.400 74.800 ;
        RECT 225.400 74.200 275.600 74.400 ;
        RECT 24.400 73.800 74.400 74.200 ;
        RECT 24.200 73.600 74.400 73.800 ;
        RECT 225.600 73.800 275.600 74.200 ;
        RECT 225.600 73.600 275.800 73.800 ;
        RECT 24.200 73.200 74.200 73.600 ;
        RECT 24.000 73.000 74.200 73.200 ;
        RECT 225.800 73.200 275.800 73.600 ;
        RECT 225.800 73.000 276.000 73.200 ;
        RECT 24.000 72.600 74.000 73.000 ;
        RECT 23.800 72.400 74.000 72.600 ;
        RECT 226.000 72.600 276.000 73.000 ;
        RECT 226.000 72.400 276.200 72.600 ;
        RECT 23.800 72.000 73.800 72.400 ;
        RECT 23.500 71.800 73.800 72.000 ;
        RECT 226.200 72.000 276.200 72.400 ;
        RECT 226.200 71.800 276.500 72.000 ;
        RECT 23.500 71.400 73.500 71.800 ;
        RECT 23.300 71.200 73.500 71.400 ;
        RECT 226.500 71.400 276.500 71.800 ;
        RECT 226.500 71.200 276.700 71.400 ;
        RECT 23.300 70.800 73.300 71.200 ;
        RECT 23.100 70.600 73.300 70.800 ;
        RECT 226.700 70.800 276.700 71.200 ;
        RECT 226.700 70.600 276.900 70.800 ;
        RECT 23.100 70.200 73.100 70.600 ;
        RECT 22.800 70.000 73.100 70.200 ;
        RECT 226.900 70.200 276.900 70.600 ;
        RECT 226.900 70.000 277.200 70.200 ;
        RECT 22.800 69.600 72.800 70.000 ;
        RECT 22.600 69.400 72.800 69.600 ;
        RECT 227.200 69.600 277.200 70.000 ;
        RECT 227.200 69.400 277.400 69.600 ;
        RECT 22.600 69.000 72.600 69.400 ;
        RECT 22.400 68.800 72.600 69.000 ;
        RECT 227.400 69.000 277.400 69.400 ;
        RECT 227.400 68.800 277.600 69.000 ;
        RECT 22.400 68.400 72.400 68.800 ;
        RECT 22.200 68.200 72.400 68.400 ;
        RECT 227.600 68.400 277.600 68.800 ;
        RECT 227.600 68.200 277.800 68.400 ;
        RECT 22.200 67.800 72.200 68.200 ;
        RECT 22.000 67.600 72.200 67.800 ;
        RECT 227.800 67.800 277.800 68.200 ;
        RECT 227.800 67.600 278.000 67.800 ;
        RECT 22.000 67.200 72.000 67.600 ;
        RECT 21.700 67.000 72.000 67.200 ;
        RECT 228.000 67.200 278.000 67.600 ;
        RECT 228.000 67.000 278.300 67.200 ;
        RECT 21.700 66.600 71.700 67.000 ;
        RECT 21.500 66.400 71.700 66.600 ;
        RECT 228.300 66.600 278.300 67.000 ;
        RECT 228.300 66.400 278.500 66.600 ;
        RECT 21.500 66.000 71.500 66.400 ;
        RECT 21.300 65.800 71.500 66.000 ;
        RECT 228.500 66.000 278.500 66.400 ;
        RECT 228.500 65.800 278.700 66.000 ;
        RECT 21.300 65.400 71.300 65.800 ;
        RECT 21.000 65.200 71.300 65.400 ;
        RECT 228.700 65.400 278.700 65.800 ;
        RECT 228.700 65.200 279.000 65.400 ;
        RECT 21.000 64.800 71.000 65.200 ;
        RECT 20.800 64.600 71.000 64.800 ;
        RECT 229.000 64.800 279.000 65.200 ;
        RECT 229.000 64.600 279.200 64.800 ;
        RECT 20.800 64.200 70.800 64.600 ;
        RECT 20.600 64.000 70.800 64.200 ;
        RECT 229.200 64.200 279.200 64.600 ;
        RECT 229.200 64.000 279.400 64.200 ;
        RECT 20.600 63.600 70.600 64.000 ;
        RECT 20.400 63.400 70.600 63.600 ;
        RECT 229.400 63.600 279.400 64.000 ;
        RECT 229.400 63.400 279.600 63.600 ;
        RECT 20.400 63.000 70.400 63.400 ;
        RECT 20.100 62.800 70.400 63.000 ;
        RECT 229.600 63.000 279.600 63.400 ;
        RECT 229.600 62.800 279.800 63.000 ;
        RECT 20.100 62.400 70.100 62.800 ;
        RECT 19.900 62.200 70.100 62.400 ;
        RECT 229.900 62.400 279.800 62.800 ;
        RECT 229.900 62.200 280.100 62.400 ;
        RECT 19.900 61.800 69.900 62.200 ;
        RECT 19.700 61.600 69.900 61.800 ;
        RECT 230.100 61.800 280.100 62.200 ;
        RECT 230.100 61.600 280.300 61.800 ;
        RECT 19.700 61.200 69.700 61.600 ;
        RECT 19.500 61.000 69.700 61.200 ;
        RECT 230.300 61.200 280.300 61.600 ;
        RECT 230.300 61.000 280.500 61.200 ;
        RECT 19.500 60.600 69.500 61.000 ;
        RECT 19.200 60.400 69.500 60.600 ;
        RECT 230.500 60.600 280.500 61.000 ;
        RECT 230.500 60.400 280.800 60.600 ;
        RECT 19.200 60.000 69.200 60.400 ;
        RECT 19.000 59.800 69.200 60.000 ;
        RECT 230.800 60.000 280.800 60.400 ;
        RECT 230.800 59.800 281.000 60.000 ;
        RECT 19.000 59.400 69.000 59.800 ;
        RECT 18.800 59.200 69.000 59.400 ;
        RECT 231.000 59.400 281.000 59.800 ;
        RECT 231.000 59.200 281.200 59.400 ;
        RECT 18.800 58.800 68.800 59.200 ;
        RECT 18.600 58.600 68.800 58.800 ;
        RECT 231.200 58.800 281.200 59.200 ;
        RECT 231.200 58.600 281.400 58.800 ;
        RECT 18.600 58.200 68.600 58.600 ;
        RECT 18.300 58.000 68.600 58.200 ;
        RECT 231.400 58.200 281.400 58.600 ;
        RECT 231.400 58.000 281.600 58.200 ;
        RECT 18.300 57.600 68.400 58.000 ;
        RECT 18.100 57.400 68.400 57.600 ;
        RECT 231.600 57.600 281.600 58.000 ;
        RECT 231.600 57.400 281.900 57.600 ;
        RECT 18.100 57.000 68.100 57.400 ;
        RECT 17.900 56.800 68.100 57.000 ;
        RECT 231.900 57.000 281.900 57.400 ;
        RECT 231.900 56.800 282.100 57.000 ;
        RECT 17.900 56.400 67.900 56.800 ;
        RECT 17.700 56.200 67.900 56.400 ;
        RECT 232.100 56.400 282.100 56.800 ;
        RECT 232.100 56.200 282.300 56.400 ;
        RECT 17.700 55.800 67.700 56.200 ;
        RECT 17.500 55.600 67.700 55.800 ;
        RECT 232.300 55.800 282.300 56.200 ;
        RECT 232.300 55.600 282.600 55.800 ;
        RECT 17.500 55.200 67.400 55.600 ;
        RECT 17.200 55.000 67.400 55.200 ;
        RECT 232.600 55.200 282.600 55.600 ;
        RECT 232.600 55.000 282.800 55.200 ;
        RECT 17.200 54.600 67.200 55.000 ;
        RECT 17.000 54.400 67.200 54.600 ;
        RECT 232.800 54.600 282.800 55.000 ;
        RECT 232.800 54.400 283.000 54.600 ;
        RECT 17.000 54.000 67.000 54.400 ;
        RECT 16.800 53.800 67.000 54.000 ;
        RECT 233.000 54.000 283.000 54.400 ;
        RECT 233.000 53.800 283.200 54.000 ;
        RECT 16.800 53.400 66.800 53.800 ;
        RECT 16.500 53.200 66.800 53.400 ;
        RECT 233.200 53.400 283.200 53.800 ;
        RECT 233.200 53.200 283.400 53.400 ;
        RECT 16.500 52.800 66.600 53.200 ;
        RECT 16.300 52.600 66.600 52.800 ;
        RECT 233.400 52.800 283.400 53.200 ;
        RECT 233.400 52.600 283.700 52.800 ;
        RECT 16.300 52.200 66.300 52.600 ;
        RECT 16.100 52.000 66.300 52.200 ;
        RECT 233.700 52.200 283.700 52.600 ;
        RECT 233.700 52.000 283.900 52.200 ;
        RECT 16.100 51.600 66.100 52.000 ;
        RECT 15.900 51.400 66.100 51.600 ;
        RECT 233.900 51.600 283.900 52.000 ;
        RECT 233.900 51.400 284.100 51.600 ;
        RECT 15.900 51.000 65.900 51.400 ;
        RECT 15.600 50.800 65.900 51.000 ;
        RECT 234.100 51.000 284.100 51.400 ;
        RECT 234.100 50.800 284.400 51.000 ;
        RECT 15.600 50.400 65.600 50.800 ;
        RECT 15.400 50.200 65.600 50.400 ;
        RECT 234.400 50.400 284.400 50.800 ;
        RECT 234.400 50.200 284.600 50.400 ;
        RECT 15.400 49.800 65.400 50.200 ;
        RECT 15.200 49.600 65.400 49.800 ;
        RECT 234.600 49.800 284.600 50.200 ;
        RECT 234.600 49.600 284.800 49.800 ;
        RECT 15.200 49.200 65.200 49.600 ;
        RECT 15.000 49.000 65.200 49.200 ;
        RECT 234.800 49.200 284.800 49.600 ;
        RECT 234.800 49.000 285.000 49.200 ;
        RECT 15.000 48.600 65.000 49.000 ;
        RECT 14.800 48.400 65.000 48.600 ;
        RECT 235.000 48.600 285.000 49.000 ;
        RECT 235.000 48.400 285.200 48.600 ;
        RECT 14.800 48.000 64.800 48.400 ;
        RECT 14.500 47.800 64.800 48.000 ;
        RECT 235.200 48.000 285.200 48.400 ;
        RECT 235.200 47.800 285.500 48.000 ;
        RECT 14.500 47.400 64.500 47.800 ;
        RECT 14.300 47.200 64.500 47.400 ;
        RECT 235.500 47.400 285.500 47.800 ;
        RECT 235.500 47.200 285.700 47.400 ;
        RECT 14.300 46.800 64.300 47.200 ;
        RECT 14.100 46.600 64.300 46.800 ;
        RECT 235.700 46.800 285.700 47.200 ;
        RECT 235.700 46.600 285.900 46.800 ;
        RECT 14.100 46.200 64.100 46.600 ;
        RECT 13.800 46.000 64.100 46.200 ;
        RECT 235.900 46.200 285.900 46.600 ;
        RECT 235.900 46.000 286.200 46.200 ;
        RECT 13.800 45.600 63.800 46.000 ;
        RECT 13.600 45.400 63.800 45.600 ;
        RECT 236.100 45.600 286.200 46.000 ;
        RECT 236.100 45.400 286.400 45.600 ;
        RECT 13.600 45.000 63.600 45.400 ;
        RECT 13.400 44.800 63.600 45.000 ;
        RECT 236.400 45.000 286.400 45.400 ;
        RECT 236.400 44.800 286.600 45.000 ;
        RECT 13.400 44.400 63.400 44.800 ;
        RECT 13.200 44.200 63.400 44.400 ;
        RECT 236.600 44.400 286.600 44.800 ;
        RECT 236.600 44.200 286.800 44.400 ;
        RECT 13.200 43.800 63.200 44.200 ;
        RECT 13.000 43.600 63.200 43.800 ;
        RECT 236.800 43.800 286.800 44.200 ;
        RECT 236.800 43.600 287.000 43.800 ;
        RECT 13.000 43.200 63.000 43.600 ;
        RECT 12.700 43.000 63.000 43.200 ;
        RECT 237.000 43.200 287.000 43.600 ;
        RECT 237.000 43.000 287.300 43.200 ;
        RECT 12.700 42.600 62.700 43.000 ;
        RECT 12.500 42.400 62.700 42.600 ;
        RECT 237.300 42.600 287.300 43.000 ;
        RECT 237.300 42.400 287.500 42.600 ;
        RECT 12.500 42.000 62.500 42.400 ;
        RECT 12.300 41.800 62.500 42.000 ;
        RECT 237.500 42.000 287.500 42.400 ;
        RECT 237.500 41.800 287.700 42.000 ;
        RECT 12.300 41.400 62.300 41.800 ;
        RECT 12.000 41.200 62.300 41.400 ;
        RECT 237.700 41.400 287.700 41.800 ;
        RECT 237.700 41.200 288.000 41.400 ;
        RECT 12.000 40.800 62.000 41.200 ;
        RECT 11.800 40.600 62.000 40.800 ;
        RECT 238.000 40.800 288.000 41.200 ;
        RECT 238.000 40.600 288.200 40.800 ;
        RECT 11.800 40.200 61.800 40.600 ;
        RECT 11.600 40.000 61.800 40.200 ;
        RECT 238.200 40.200 288.200 40.600 ;
        RECT 238.200 40.000 288.400 40.200 ;
        RECT 11.600 39.600 61.600 40.000 ;
        RECT 11.400 39.400 61.600 39.600 ;
        RECT 238.400 39.600 288.400 40.000 ;
        RECT 238.400 39.400 288.600 39.600 ;
        RECT 11.400 39.000 61.400 39.400 ;
        RECT 11.100 38.800 61.400 39.000 ;
        RECT 238.600 39.000 288.600 39.400 ;
        RECT 238.600 38.800 288.800 39.000 ;
        RECT 11.100 38.400 61.100 38.800 ;
        RECT 10.900 38.200 61.100 38.400 ;
        RECT 238.900 38.400 288.800 38.800 ;
        RECT 238.900 38.200 289.100 38.400 ;
        RECT 10.900 37.800 60.900 38.200 ;
        RECT 10.700 37.600 60.900 37.800 ;
        RECT 239.100 37.800 289.100 38.200 ;
        RECT 239.100 37.600 289.300 37.800 ;
        RECT 10.700 37.200 60.700 37.600 ;
        RECT 10.500 37.000 60.700 37.200 ;
        RECT 239.300 37.200 289.300 37.600 ;
        RECT 239.300 37.000 289.500 37.200 ;
        RECT 10.500 36.600 60.500 37.000 ;
        RECT 10.200 36.400 60.500 36.600 ;
        RECT 239.500 36.600 289.500 37.000 ;
        RECT 239.500 36.400 289.800 36.600 ;
        RECT 10.200 36.000 60.200 36.400 ;
        RECT 10.000 35.800 60.200 36.000 ;
        RECT 239.800 36.000 289.800 36.400 ;
        RECT 239.800 35.800 290.000 36.000 ;
        RECT 10.000 35.400 60.000 35.800 ;
        RECT 9.800 35.200 60.000 35.400 ;
        RECT 240.000 35.400 290.000 35.800 ;
        RECT 240.000 35.200 290.200 35.400 ;
        RECT 9.800 34.800 59.800 35.200 ;
        RECT 9.600 34.600 59.800 34.800 ;
        RECT 240.200 34.800 290.200 35.200 ;
        RECT 240.200 34.600 290.400 34.800 ;
        RECT 9.600 34.200 59.600 34.600 ;
        RECT 9.300 34.000 59.600 34.200 ;
        RECT 240.400 34.200 290.400 34.600 ;
        RECT 240.400 34.000 290.600 34.200 ;
        RECT 9.300 33.600 59.300 34.000 ;
        RECT 9.100 33.400 59.300 33.600 ;
        RECT 240.600 33.600 290.600 34.000 ;
        RECT 240.600 33.400 290.900 33.600 ;
        RECT 9.100 33.000 59.100 33.400 ;
        RECT 8.900 32.800 59.100 33.000 ;
        RECT 240.900 33.000 290.900 33.400 ;
        RECT 240.900 32.800 291.100 33.000 ;
        RECT 8.900 32.400 58.900 32.800 ;
        RECT 8.700 32.200 58.900 32.400 ;
        RECT 241.100 32.400 291.100 32.800 ;
        RECT 241.100 32.200 291.300 32.400 ;
        RECT 8.700 31.800 58.700 32.200 ;
        RECT 8.500 31.600 58.700 31.800 ;
        RECT 241.300 31.800 291.300 32.200 ;
        RECT 241.300 31.600 291.600 31.800 ;
        RECT 8.500 31.200 58.400 31.600 ;
        RECT 8.200 31.000 58.400 31.200 ;
        RECT 241.600 31.200 291.600 31.600 ;
        RECT 241.600 31.000 291.800 31.200 ;
        RECT 8.200 30.600 58.200 31.000 ;
        RECT 8.000 30.400 58.200 30.600 ;
        RECT 241.800 30.600 291.800 31.000 ;
        RECT 241.800 30.400 292.000 30.600 ;
        RECT 8.000 30.000 58.000 30.400 ;
        RECT 7.800 29.800 58.000 30.000 ;
        RECT 242.000 30.000 292.000 30.400 ;
        RECT 242.000 29.800 292.200 30.000 ;
        RECT 7.800 29.400 57.800 29.800 ;
        RECT 7.500 29.200 57.800 29.400 ;
        RECT 242.200 29.400 292.200 29.800 ;
        RECT 242.200 29.200 292.400 29.400 ;
        RECT 7.500 28.800 57.600 29.200 ;
        RECT 7.300 28.600 57.600 28.800 ;
        RECT 242.400 28.800 292.400 29.200 ;
        RECT 242.400 28.600 292.700 28.800 ;
        RECT 7.300 28.200 57.300 28.600 ;
        RECT 7.100 28.000 57.300 28.200 ;
        RECT 242.700 28.200 292.700 28.600 ;
        RECT 242.700 28.000 292.900 28.200 ;
        RECT 7.100 27.600 57.100 28.000 ;
        RECT 6.900 27.400 57.100 27.600 ;
        RECT 242.900 27.600 292.900 28.000 ;
        RECT 242.900 27.400 293.100 27.600 ;
        RECT 6.900 27.000 56.900 27.400 ;
        RECT 6.600 26.800 56.900 27.000 ;
        RECT 243.100 27.000 293.100 27.400 ;
        RECT 243.100 26.800 293.400 27.000 ;
        RECT 6.600 26.400 56.600 26.800 ;
        RECT 6.400 26.200 56.600 26.400 ;
        RECT 243.400 26.400 293.400 26.800 ;
        RECT 243.400 26.200 293.600 26.400 ;
        RECT 6.400 25.800 56.400 26.200 ;
        RECT 6.200 25.600 56.400 25.800 ;
        RECT 243.600 25.800 293.600 26.200 ;
        RECT 243.600 25.600 293.800 25.800 ;
        RECT 6.200 25.200 56.200 25.600 ;
        RECT 6.000 25.000 56.200 25.200 ;
        RECT 243.800 25.200 293.800 25.600 ;
        RECT 243.800 25.000 294.000 25.200 ;
        RECT 6.000 24.600 56.000 25.000 ;
        RECT 5.800 24.400 56.000 24.600 ;
        RECT 244.000 24.600 294.000 25.000 ;
        RECT 244.000 24.400 294.200 24.600 ;
        RECT 5.800 24.000 55.800 24.400 ;
        RECT 5.500 23.800 55.800 24.000 ;
        RECT 244.200 24.000 294.200 24.400 ;
        RECT 244.200 23.800 294.500 24.000 ;
        RECT 5.500 23.400 55.500 23.800 ;
        RECT 5.300 23.200 55.500 23.400 ;
        RECT 244.500 23.400 294.500 23.800 ;
        RECT 244.500 23.200 294.700 23.400 ;
        RECT 5.300 22.800 55.300 23.200 ;
        RECT 5.100 22.600 55.300 22.800 ;
        RECT 244.700 22.800 294.700 23.200 ;
        RECT 244.700 22.600 294.900 22.800 ;
        RECT 5.100 22.200 55.100 22.600 ;
        RECT 4.800 22.000 55.100 22.200 ;
        RECT 244.900 22.200 294.900 22.600 ;
        RECT 244.900 22.000 295.200 22.200 ;
        RECT 4.800 21.600 54.800 22.000 ;
        RECT 4.600 21.400 54.800 21.600 ;
        RECT 245.100 21.600 295.200 22.000 ;
        RECT 245.100 21.400 295.400 21.600 ;
        RECT 4.600 21.000 54.600 21.400 ;
        RECT 4.400 20.800 54.600 21.000 ;
        RECT 245.400 21.000 295.400 21.400 ;
        RECT 245.400 20.800 295.600 21.000 ;
        RECT 4.400 20.400 54.400 20.800 ;
        RECT 4.200 20.200 54.400 20.400 ;
        RECT 245.600 20.400 295.600 20.800 ;
        RECT 245.600 20.200 295.800 20.400 ;
        RECT 4.200 19.800 54.200 20.200 ;
        RECT 4.000 19.600 54.200 19.800 ;
        RECT 245.800 19.800 295.800 20.200 ;
        RECT 245.800 19.600 296.000 19.800 ;
        RECT 4.000 19.200 54.000 19.600 ;
        RECT 3.700 19.000 54.000 19.200 ;
        RECT 246.000 19.200 296.000 19.600 ;
        RECT 246.000 19.000 296.300 19.200 ;
        RECT 3.700 18.600 53.700 19.000 ;
        RECT 3.500 18.400 53.700 18.600 ;
        RECT 246.300 18.600 296.300 19.000 ;
        RECT 246.300 18.400 296.500 18.600 ;
        RECT 3.500 18.000 53.500 18.400 ;
        RECT 3.300 17.800 53.500 18.000 ;
        RECT 246.500 18.000 296.500 18.400 ;
        RECT 246.500 17.800 296.700 18.000 ;
        RECT 3.300 17.400 53.300 17.800 ;
        RECT 3.000 17.200 53.300 17.400 ;
        RECT 246.700 17.400 296.700 17.800 ;
        RECT 246.700 17.200 297.000 17.400 ;
        RECT 3.000 16.800 53.000 17.200 ;
        RECT 2.800 16.600 53.000 16.800 ;
        RECT 247.000 16.800 297.000 17.200 ;
        RECT 247.000 16.600 297.200 16.800 ;
        RECT 2.800 16.200 52.800 16.600 ;
        RECT 2.600 16.000 52.800 16.200 ;
        RECT 247.200 16.200 297.200 16.600 ;
        RECT 247.200 16.000 297.400 16.200 ;
        RECT 2.600 15.600 52.600 16.000 ;
        RECT 2.400 15.400 52.600 15.600 ;
        RECT 247.400 15.600 297.400 16.000 ;
        RECT 247.400 15.400 297.600 15.600 ;
        RECT 2.400 15.000 52.400 15.400 ;
        RECT 2.100 14.800 52.400 15.000 ;
        RECT 247.600 15.000 297.600 15.400 ;
        RECT 247.600 14.800 297.800 15.000 ;
        RECT 2.100 14.400 52.100 14.800 ;
        RECT 1.900 14.200 52.100 14.400 ;
        RECT 247.900 14.400 297.800 14.800 ;
        RECT 247.900 14.200 298.100 14.400 ;
        RECT 1.900 13.800 51.900 14.200 ;
        RECT 1.700 13.600 51.900 13.800 ;
        RECT 248.100 13.800 298.100 14.200 ;
        RECT 248.100 13.600 298.300 13.800 ;
        RECT 1.700 13.200 51.700 13.600 ;
        RECT 1.500 13.000 51.700 13.200 ;
        RECT 248.300 13.200 298.300 13.600 ;
        RECT 248.300 13.000 298.500 13.200 ;
        RECT 1.500 12.400 51.500 13.000 ;
        RECT 248.500 12.400 298.500 13.000 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER Metal5 ;
        RECT 337.500 342.600 342.500 344.700 ;
        RECT 315.000 342.000 365.000 342.600 ;
        RECT 315.000 341.400 365.400 342.000 ;
        RECT 315.000 340.800 365.800 341.400 ;
        RECT 315.000 340.200 366.200 340.800 ;
        RECT 315.000 339.600 366.600 340.200 ;
        RECT 315.000 339.000 367.000 339.600 ;
        RECT 315.000 338.400 367.400 339.000 ;
        RECT 315.000 337.800 367.800 338.400 ;
        RECT 315.000 337.200 368.200 337.800 ;
        RECT 315.000 336.600 368.600 337.200 ;
        RECT 315.000 336.000 369.000 336.600 ;
        RECT 315.000 335.400 369.400 336.000 ;
        RECT 315.000 334.800 369.800 335.400 ;
        RECT 315.000 334.200 370.200 334.800 ;
        RECT 315.000 333.600 370.600 334.200 ;
        RECT 315.000 333.000 371.000 333.600 ;
        RECT 315.000 332.400 371.400 333.000 ;
        RECT 315.000 331.800 371.800 332.400 ;
        RECT 315.000 331.200 372.200 331.800 ;
        RECT 315.000 330.600 372.600 331.200 ;
        RECT 315.000 330.000 373.000 330.600 ;
        RECT 315.000 329.400 373.400 330.000 ;
        RECT 315.000 328.800 373.800 329.400 ;
        RECT 315.000 328.200 374.200 328.800 ;
        RECT 315.000 327.600 374.600 328.200 ;
        RECT 315.000 327.000 375.000 327.600 ;
        RECT 315.000 326.400 375.400 327.000 ;
        RECT 315.000 325.800 375.800 326.400 ;
        RECT 315.000 325.200 376.200 325.800 ;
        RECT 315.000 324.600 376.600 325.200 ;
        RECT 315.000 324.000 377.000 324.600 ;
        RECT 315.000 323.400 377.400 324.000 ;
        RECT 315.000 322.800 377.800 323.400 ;
        RECT 315.000 322.200 378.200 322.800 ;
        RECT 315.000 321.600 378.600 322.200 ;
        RECT 315.000 321.000 379.000 321.600 ;
        RECT 315.000 320.400 379.400 321.000 ;
        RECT 315.000 319.800 379.800 320.400 ;
        RECT 315.000 319.200 380.200 319.800 ;
        RECT 315.000 318.600 380.600 319.200 ;
        RECT 315.000 318.000 381.000 318.600 ;
        RECT 315.000 317.400 381.400 318.000 ;
        RECT 315.000 316.800 381.800 317.400 ;
        RECT 315.000 316.200 382.200 316.800 ;
        RECT 315.000 315.600 382.600 316.200 ;
        RECT 315.000 315.000 383.000 315.600 ;
        RECT 315.000 314.400 383.400 315.000 ;
        RECT 315.000 313.800 383.800 314.400 ;
        RECT 315.000 313.200 384.200 313.800 ;
        RECT 315.000 312.600 384.600 313.200 ;
        RECT 315.000 312.000 385.000 312.600 ;
        RECT 315.000 311.400 385.400 312.000 ;
        RECT 315.000 310.800 385.800 311.400 ;
        RECT 315.000 310.200 386.200 310.800 ;
        RECT 315.000 309.600 386.600 310.200 ;
        RECT 315.000 309.000 387.000 309.600 ;
        RECT 315.000 308.400 387.400 309.000 ;
        RECT 315.000 307.800 387.800 308.400 ;
        RECT 315.000 307.200 388.200 307.800 ;
        RECT 315.000 306.600 388.600 307.200 ;
        RECT 315.000 306.000 389.000 306.600 ;
        RECT 315.000 305.400 389.400 306.000 ;
        RECT 315.000 304.800 389.800 305.400 ;
        RECT 315.000 304.200 390.200 304.800 ;
        RECT 315.000 303.600 390.600 304.200 ;
        RECT 315.000 303.000 391.000 303.600 ;
        RECT 315.000 302.400 391.400 303.000 ;
        RECT 315.000 301.800 391.800 302.400 ;
        RECT 315.000 301.200 392.200 301.800 ;
        RECT 315.000 300.600 392.600 301.200 ;
        RECT 315.000 300.000 393.000 300.600 ;
        RECT 315.000 299.400 393.400 300.000 ;
        RECT 315.000 298.800 393.800 299.400 ;
        RECT 315.000 298.200 394.200 298.800 ;
        RECT 315.000 297.600 394.600 298.200 ;
        RECT 315.000 297.000 395.000 297.600 ;
        RECT 315.000 296.400 395.400 297.000 ;
        RECT 315.000 295.800 395.800 296.400 ;
        RECT 315.000 295.200 396.200 295.800 ;
        RECT 315.000 294.600 396.600 295.200 ;
        RECT 315.000 294.000 397.000 294.600 ;
        RECT 315.000 293.400 397.400 294.000 ;
        RECT 315.000 292.800 397.800 293.400 ;
        RECT 315.000 292.200 398.200 292.800 ;
        RECT 315.000 291.600 398.600 292.200 ;
        RECT 315.000 291.000 399.000 291.600 ;
        RECT 315.000 290.400 399.400 291.000 ;
        RECT 315.000 289.800 399.800 290.400 ;
        RECT 315.000 289.200 400.200 289.800 ;
        RECT 315.000 288.600 400.600 289.200 ;
        RECT 315.000 288.000 401.000 288.600 ;
        RECT 315.000 287.400 401.400 288.000 ;
        RECT 315.000 286.800 401.800 287.400 ;
        RECT 315.000 286.200 402.200 286.800 ;
        RECT 315.000 285.600 402.600 286.200 ;
        RECT 315.000 285.000 403.000 285.600 ;
        RECT 315.000 284.400 403.400 285.000 ;
        RECT 315.000 283.800 403.800 284.400 ;
        RECT 315.000 283.200 404.200 283.800 ;
        RECT 315.000 282.600 404.600 283.200 ;
        RECT 315.000 282.000 405.000 282.600 ;
        RECT 315.000 281.400 405.400 282.000 ;
        RECT 315.000 280.800 405.800 281.400 ;
        RECT 315.000 280.200 406.200 280.800 ;
        RECT 315.000 279.600 406.600 280.200 ;
        RECT 315.000 279.000 407.000 279.600 ;
        RECT 315.000 278.400 407.400 279.000 ;
        RECT 315.000 277.800 407.800 278.400 ;
        RECT 315.000 277.200 408.200 277.800 ;
        RECT 315.000 276.600 408.600 277.200 ;
        RECT 315.000 276.000 409.000 276.600 ;
        RECT 315.000 275.400 409.400 276.000 ;
        RECT 315.000 274.800 409.800 275.400 ;
        RECT 315.000 274.200 410.200 274.800 ;
        RECT 315.000 273.600 410.600 274.200 ;
        RECT 315.000 273.000 411.000 273.600 ;
        RECT 315.000 272.400 411.400 273.000 ;
        RECT 315.000 271.800 411.800 272.400 ;
        RECT 315.000 271.200 412.200 271.800 ;
        RECT 315.000 270.600 412.600 271.200 ;
        RECT 315.000 270.000 413.000 270.600 ;
        RECT 315.000 269.400 413.400 270.000 ;
        RECT 315.000 268.800 413.800 269.400 ;
        RECT 315.000 268.200 414.200 268.800 ;
        RECT 315.000 267.600 414.600 268.200 ;
        RECT 315.000 267.000 415.000 267.600 ;
        RECT 315.000 266.800 415.400 267.000 ;
        RECT 315.000 12.400 365.000 266.800 ;
        RECT 365.400 266.400 415.400 266.800 ;
        RECT 365.400 266.200 415.800 266.400 ;
        RECT 365.800 265.800 415.800 266.200 ;
        RECT 365.800 265.600 416.200 265.800 ;
        RECT 366.200 265.200 416.200 265.600 ;
        RECT 366.200 265.000 416.600 265.200 ;
        RECT 366.600 264.600 416.600 265.000 ;
        RECT 366.600 264.400 417.000 264.600 ;
        RECT 367.000 264.000 417.000 264.400 ;
        RECT 367.000 263.800 417.400 264.000 ;
        RECT 367.400 263.400 417.400 263.800 ;
        RECT 367.400 263.200 417.800 263.400 ;
        RECT 367.800 262.800 417.800 263.200 ;
        RECT 367.800 262.600 418.200 262.800 ;
        RECT 368.200 262.200 418.200 262.600 ;
        RECT 368.200 262.000 418.600 262.200 ;
        RECT 368.600 261.600 418.600 262.000 ;
        RECT 368.600 261.400 419.000 261.600 ;
        RECT 369.000 261.000 419.000 261.400 ;
        RECT 369.000 260.800 419.400 261.000 ;
        RECT 369.400 260.400 419.400 260.800 ;
        RECT 369.400 260.200 419.800 260.400 ;
        RECT 369.800 259.800 419.800 260.200 ;
        RECT 369.800 259.600 420.200 259.800 ;
        RECT 370.200 259.200 420.200 259.600 ;
        RECT 370.200 259.000 420.600 259.200 ;
        RECT 370.600 258.600 420.600 259.000 ;
        RECT 370.600 258.400 421.000 258.600 ;
        RECT 371.000 258.000 421.000 258.400 ;
        RECT 371.000 257.800 421.400 258.000 ;
        RECT 371.400 257.400 421.400 257.800 ;
        RECT 371.400 257.200 421.800 257.400 ;
        RECT 371.800 256.800 421.800 257.200 ;
        RECT 371.800 256.600 422.200 256.800 ;
        RECT 372.200 256.200 422.200 256.600 ;
        RECT 372.200 256.000 422.600 256.200 ;
        RECT 372.600 255.600 422.600 256.000 ;
        RECT 372.600 255.400 423.000 255.600 ;
        RECT 373.000 255.000 423.000 255.400 ;
        RECT 373.000 254.800 423.400 255.000 ;
        RECT 373.400 254.400 423.400 254.800 ;
        RECT 373.400 254.200 423.800 254.400 ;
        RECT 373.800 253.800 423.800 254.200 ;
        RECT 373.800 253.600 424.200 253.800 ;
        RECT 374.200 253.200 424.200 253.600 ;
        RECT 374.200 253.000 424.600 253.200 ;
        RECT 374.600 252.600 424.600 253.000 ;
        RECT 374.600 252.400 425.000 252.600 ;
        RECT 375.000 252.000 425.000 252.400 ;
        RECT 375.000 251.800 425.400 252.000 ;
        RECT 375.400 251.400 425.400 251.800 ;
        RECT 375.400 251.200 425.800 251.400 ;
        RECT 375.800 250.800 425.800 251.200 ;
        RECT 375.800 250.600 426.200 250.800 ;
        RECT 376.200 250.200 426.200 250.600 ;
        RECT 376.200 250.000 426.600 250.200 ;
        RECT 376.600 249.600 426.600 250.000 ;
        RECT 376.600 249.400 427.000 249.600 ;
        RECT 377.000 249.000 427.000 249.400 ;
        RECT 377.000 248.800 427.400 249.000 ;
        RECT 377.400 248.400 427.400 248.800 ;
        RECT 377.400 248.200 427.800 248.400 ;
        RECT 377.800 247.800 427.800 248.200 ;
        RECT 377.800 247.600 428.200 247.800 ;
        RECT 378.200 247.200 428.200 247.600 ;
        RECT 378.200 247.000 428.600 247.200 ;
        RECT 378.600 246.600 428.600 247.000 ;
        RECT 378.600 246.400 429.000 246.600 ;
        RECT 379.000 246.000 429.000 246.400 ;
        RECT 379.000 245.800 429.400 246.000 ;
        RECT 379.400 245.400 429.400 245.800 ;
        RECT 379.400 245.200 429.800 245.400 ;
        RECT 379.800 244.800 429.800 245.200 ;
        RECT 379.800 244.600 430.200 244.800 ;
        RECT 380.200 244.200 430.200 244.600 ;
        RECT 380.200 244.000 430.600 244.200 ;
        RECT 380.600 243.600 430.600 244.000 ;
        RECT 380.600 243.400 431.000 243.600 ;
        RECT 381.000 243.000 431.000 243.400 ;
        RECT 381.000 242.800 431.400 243.000 ;
        RECT 381.400 242.400 431.400 242.800 ;
        RECT 381.400 242.200 431.800 242.400 ;
        RECT 381.800 241.800 431.800 242.200 ;
        RECT 381.800 241.600 432.200 241.800 ;
        RECT 382.200 241.200 432.200 241.600 ;
        RECT 382.200 241.000 432.600 241.200 ;
        RECT 382.600 240.600 432.600 241.000 ;
        RECT 382.600 240.400 433.000 240.600 ;
        RECT 383.000 240.000 433.000 240.400 ;
        RECT 383.000 239.800 433.400 240.000 ;
        RECT 383.400 239.400 433.400 239.800 ;
        RECT 383.400 239.200 433.800 239.400 ;
        RECT 383.800 238.800 433.800 239.200 ;
        RECT 383.800 238.600 434.200 238.800 ;
        RECT 384.200 238.200 434.200 238.600 ;
        RECT 384.200 238.000 434.600 238.200 ;
        RECT 384.600 237.600 434.600 238.000 ;
        RECT 384.600 237.400 435.000 237.600 ;
        RECT 385.000 237.000 435.000 237.400 ;
        RECT 385.000 236.800 435.400 237.000 ;
        RECT 385.400 236.400 435.400 236.800 ;
        RECT 385.400 236.200 435.800 236.400 ;
        RECT 385.800 235.800 435.800 236.200 ;
        RECT 385.800 235.600 436.200 235.800 ;
        RECT 386.200 235.200 436.200 235.600 ;
        RECT 386.200 235.000 436.600 235.200 ;
        RECT 386.600 234.600 436.600 235.000 ;
        RECT 386.600 234.400 437.000 234.600 ;
        RECT 387.000 234.000 437.000 234.400 ;
        RECT 387.000 233.800 437.400 234.000 ;
        RECT 387.400 233.400 437.400 233.800 ;
        RECT 387.400 233.200 437.800 233.400 ;
        RECT 387.800 232.800 437.800 233.200 ;
        RECT 387.800 232.600 438.200 232.800 ;
        RECT 388.200 232.200 438.200 232.600 ;
        RECT 388.200 232.000 438.600 232.200 ;
        RECT 388.600 231.600 438.600 232.000 ;
        RECT 388.600 231.400 439.000 231.600 ;
        RECT 389.000 231.000 439.000 231.400 ;
        RECT 389.000 230.800 439.400 231.000 ;
        RECT 389.400 230.400 439.400 230.800 ;
        RECT 389.400 230.200 439.800 230.400 ;
        RECT 389.800 229.800 439.800 230.200 ;
        RECT 389.800 229.600 440.200 229.800 ;
        RECT 390.200 229.200 440.200 229.600 ;
        RECT 390.200 229.000 440.600 229.200 ;
        RECT 390.600 228.600 440.600 229.000 ;
        RECT 390.600 228.400 441.000 228.600 ;
        RECT 391.000 228.000 441.000 228.400 ;
        RECT 391.000 227.800 441.400 228.000 ;
        RECT 391.400 227.400 441.400 227.800 ;
        RECT 391.400 227.200 441.800 227.400 ;
        RECT 391.800 226.800 441.800 227.200 ;
        RECT 391.800 226.600 442.200 226.800 ;
        RECT 392.200 226.200 442.200 226.600 ;
        RECT 392.200 226.000 442.600 226.200 ;
        RECT 392.600 225.600 442.600 226.000 ;
        RECT 392.600 225.400 443.000 225.600 ;
        RECT 393.000 225.000 443.000 225.400 ;
        RECT 393.000 224.800 443.400 225.000 ;
        RECT 393.400 224.400 443.400 224.800 ;
        RECT 393.400 224.200 443.800 224.400 ;
        RECT 393.800 223.800 443.800 224.200 ;
        RECT 393.800 223.600 444.200 223.800 ;
        RECT 394.200 223.200 444.200 223.600 ;
        RECT 394.200 223.000 444.600 223.200 ;
        RECT 394.600 222.600 444.600 223.000 ;
        RECT 394.600 222.400 445.000 222.600 ;
        RECT 395.000 222.000 445.000 222.400 ;
        RECT 395.000 221.800 445.400 222.000 ;
        RECT 395.400 221.400 445.400 221.800 ;
        RECT 395.400 221.200 445.800 221.400 ;
        RECT 395.800 220.800 445.800 221.200 ;
        RECT 395.800 220.600 446.200 220.800 ;
        RECT 396.200 220.200 446.200 220.600 ;
        RECT 396.200 220.000 446.600 220.200 ;
        RECT 396.600 219.600 446.600 220.000 ;
        RECT 396.600 219.400 447.000 219.600 ;
        RECT 397.000 219.000 447.000 219.400 ;
        RECT 397.000 218.800 447.400 219.000 ;
        RECT 397.400 218.400 447.400 218.800 ;
        RECT 397.400 218.200 447.800 218.400 ;
        RECT 397.800 217.800 447.800 218.200 ;
        RECT 397.800 217.600 448.200 217.800 ;
        RECT 398.200 217.200 448.200 217.600 ;
        RECT 398.200 217.000 448.600 217.200 ;
        RECT 398.600 216.600 448.600 217.000 ;
        RECT 398.600 216.400 449.000 216.600 ;
        RECT 399.000 216.000 449.000 216.400 ;
        RECT 399.000 215.800 449.400 216.000 ;
        RECT 399.400 215.400 449.400 215.800 ;
        RECT 399.400 215.200 449.800 215.400 ;
        RECT 399.800 214.800 449.800 215.200 ;
        RECT 399.800 214.600 450.200 214.800 ;
        RECT 400.200 214.200 450.200 214.600 ;
        RECT 400.200 214.000 450.600 214.200 ;
        RECT 400.600 213.600 450.600 214.000 ;
        RECT 400.600 213.400 451.000 213.600 ;
        RECT 401.000 213.000 451.000 213.400 ;
        RECT 401.000 212.800 451.400 213.000 ;
        RECT 401.400 212.400 451.400 212.800 ;
        RECT 401.400 212.200 451.800 212.400 ;
        RECT 401.800 211.800 451.800 212.200 ;
        RECT 401.800 211.600 452.200 211.800 ;
        RECT 402.200 211.200 452.200 211.600 ;
        RECT 402.200 211.000 452.600 211.200 ;
        RECT 402.600 210.600 452.600 211.000 ;
        RECT 402.600 210.400 453.000 210.600 ;
        RECT 403.000 210.000 453.000 210.400 ;
        RECT 403.000 209.800 453.400 210.000 ;
        RECT 403.400 209.400 453.400 209.800 ;
        RECT 403.400 209.200 453.800 209.400 ;
        RECT 403.800 208.800 453.800 209.200 ;
        RECT 403.800 208.600 454.200 208.800 ;
        RECT 404.200 208.200 454.200 208.600 ;
        RECT 404.200 208.000 454.600 208.200 ;
        RECT 404.600 207.600 454.600 208.000 ;
        RECT 404.600 207.400 455.000 207.600 ;
        RECT 405.000 207.000 455.000 207.400 ;
        RECT 405.000 206.800 455.400 207.000 ;
        RECT 405.400 206.400 455.400 206.800 ;
        RECT 405.400 206.200 455.800 206.400 ;
        RECT 405.800 205.800 455.800 206.200 ;
        RECT 405.800 205.600 456.200 205.800 ;
        RECT 406.200 205.200 456.200 205.600 ;
        RECT 406.200 205.000 456.600 205.200 ;
        RECT 406.600 204.600 456.600 205.000 ;
        RECT 406.600 204.400 457.000 204.600 ;
        RECT 407.000 204.000 457.000 204.400 ;
        RECT 407.000 203.800 457.400 204.000 ;
        RECT 407.400 203.400 457.400 203.800 ;
        RECT 407.400 203.200 457.800 203.400 ;
        RECT 407.800 202.800 457.800 203.200 ;
        RECT 407.800 202.600 458.200 202.800 ;
        RECT 408.200 202.200 458.200 202.600 ;
        RECT 408.200 202.000 458.600 202.200 ;
        RECT 408.600 201.600 458.600 202.000 ;
        RECT 408.600 201.400 459.000 201.600 ;
        RECT 409.000 201.000 459.000 201.400 ;
        RECT 409.000 200.800 459.400 201.000 ;
        RECT 409.400 200.400 459.400 200.800 ;
        RECT 409.400 200.200 459.800 200.400 ;
        RECT 409.800 199.800 459.800 200.200 ;
        RECT 409.800 199.600 460.200 199.800 ;
        RECT 410.200 199.200 460.200 199.600 ;
        RECT 410.200 199.000 460.600 199.200 ;
        RECT 410.600 198.600 460.600 199.000 ;
        RECT 410.600 198.400 461.000 198.600 ;
        RECT 411.000 198.000 461.000 198.400 ;
        RECT 411.000 197.800 461.400 198.000 ;
        RECT 411.400 197.400 461.400 197.800 ;
        RECT 411.400 197.200 461.800 197.400 ;
        RECT 411.800 196.800 461.800 197.200 ;
        RECT 411.800 196.600 462.200 196.800 ;
        RECT 412.200 196.200 462.200 196.600 ;
        RECT 412.200 196.000 462.600 196.200 ;
        RECT 412.600 195.600 462.600 196.000 ;
        RECT 412.600 195.400 463.000 195.600 ;
        RECT 413.000 195.000 463.000 195.400 ;
        RECT 413.000 194.800 463.400 195.000 ;
        RECT 413.400 194.400 463.400 194.800 ;
        RECT 413.400 194.200 463.800 194.400 ;
        RECT 413.800 193.800 463.800 194.200 ;
        RECT 413.800 193.600 464.200 193.800 ;
        RECT 414.200 193.200 464.200 193.600 ;
        RECT 414.200 193.000 464.600 193.200 ;
        RECT 414.600 192.600 464.600 193.000 ;
        RECT 414.600 192.400 465.000 192.600 ;
        RECT 415.000 192.000 465.000 192.400 ;
        RECT 415.000 191.800 465.400 192.000 ;
        RECT 415.400 191.400 465.400 191.800 ;
        RECT 415.400 191.200 465.800 191.400 ;
        RECT 415.800 190.800 465.800 191.200 ;
        RECT 415.800 190.600 466.200 190.800 ;
        RECT 416.200 190.200 466.200 190.600 ;
        RECT 416.200 190.000 466.600 190.200 ;
        RECT 416.600 189.600 466.600 190.000 ;
        RECT 416.600 189.400 467.000 189.600 ;
        RECT 417.000 189.000 467.000 189.400 ;
        RECT 417.000 188.800 467.400 189.000 ;
        RECT 417.400 188.400 467.400 188.800 ;
        RECT 417.400 188.200 467.800 188.400 ;
        RECT 417.800 187.800 467.800 188.200 ;
        RECT 417.800 187.600 468.200 187.800 ;
        RECT 418.200 187.200 468.200 187.600 ;
        RECT 418.200 187.000 468.600 187.200 ;
        RECT 418.600 186.600 468.600 187.000 ;
        RECT 418.600 186.400 469.000 186.600 ;
        RECT 419.000 186.000 469.000 186.400 ;
        RECT 419.000 185.800 469.400 186.000 ;
        RECT 419.400 185.400 469.400 185.800 ;
        RECT 419.400 185.200 469.800 185.400 ;
        RECT 419.800 184.800 469.800 185.200 ;
        RECT 419.800 184.600 470.200 184.800 ;
        RECT 420.200 184.200 470.200 184.600 ;
        RECT 420.200 184.000 470.600 184.200 ;
        RECT 420.600 183.600 470.600 184.000 ;
        RECT 420.600 183.400 471.000 183.600 ;
        RECT 421.000 183.000 471.000 183.400 ;
        RECT 421.000 182.800 471.400 183.000 ;
        RECT 421.400 182.400 471.400 182.800 ;
        RECT 421.400 182.200 471.800 182.400 ;
        RECT 421.800 181.800 471.800 182.200 ;
        RECT 421.800 181.600 472.200 181.800 ;
        RECT 422.200 181.200 472.200 181.600 ;
        RECT 422.200 181.000 472.600 181.200 ;
        RECT 422.600 180.600 472.600 181.000 ;
        RECT 422.600 180.400 473.000 180.600 ;
        RECT 423.000 180.000 473.000 180.400 ;
        RECT 423.000 179.800 473.400 180.000 ;
        RECT 423.400 179.400 473.400 179.800 ;
        RECT 423.400 179.200 473.800 179.400 ;
        RECT 423.800 178.800 473.800 179.200 ;
        RECT 423.800 178.600 474.200 178.800 ;
        RECT 424.200 178.200 474.200 178.600 ;
        RECT 424.200 178.000 474.600 178.200 ;
        RECT 424.600 177.600 474.600 178.000 ;
        RECT 424.600 177.400 475.000 177.600 ;
        RECT 425.000 177.000 475.000 177.400 ;
        RECT 425.000 176.800 475.400 177.000 ;
        RECT 425.400 176.400 475.400 176.800 ;
        RECT 425.400 176.200 475.800 176.400 ;
        RECT 425.800 175.800 475.800 176.200 ;
        RECT 425.800 175.600 476.200 175.800 ;
        RECT 426.200 175.200 476.200 175.600 ;
        RECT 426.200 175.000 476.600 175.200 ;
        RECT 426.600 174.600 476.600 175.000 ;
        RECT 426.600 174.400 477.000 174.600 ;
        RECT 427.000 174.000 477.000 174.400 ;
        RECT 427.000 173.800 477.400 174.000 ;
        RECT 427.400 173.400 477.400 173.800 ;
        RECT 427.400 173.200 477.800 173.400 ;
        RECT 427.800 172.800 477.800 173.200 ;
        RECT 427.800 172.600 478.200 172.800 ;
        RECT 428.200 172.200 478.200 172.600 ;
        RECT 428.200 172.000 478.600 172.200 ;
        RECT 428.600 171.600 478.600 172.000 ;
        RECT 428.600 171.400 479.000 171.600 ;
        RECT 429.000 171.000 479.000 171.400 ;
        RECT 429.000 170.800 479.400 171.000 ;
        RECT 429.400 170.400 479.400 170.800 ;
        RECT 429.400 170.200 479.800 170.400 ;
        RECT 429.800 169.800 479.800 170.200 ;
        RECT 429.800 169.600 480.200 169.800 ;
        RECT 430.200 169.200 480.200 169.600 ;
        RECT 430.200 169.000 480.600 169.200 ;
        RECT 430.600 168.600 480.600 169.000 ;
        RECT 430.600 168.400 481.000 168.600 ;
        RECT 431.000 168.000 481.000 168.400 ;
        RECT 431.000 167.800 481.400 168.000 ;
        RECT 431.400 167.400 481.400 167.800 ;
        RECT 431.400 167.200 481.800 167.400 ;
        RECT 431.800 166.800 481.800 167.200 ;
        RECT 431.800 166.600 482.200 166.800 ;
        RECT 432.200 166.200 482.200 166.600 ;
        RECT 432.200 166.000 482.600 166.200 ;
        RECT 432.600 165.600 482.600 166.000 ;
        RECT 432.600 165.400 483.000 165.600 ;
        RECT 433.000 165.000 483.000 165.400 ;
        RECT 433.000 164.800 483.400 165.000 ;
        RECT 433.400 164.400 483.400 164.800 ;
        RECT 433.400 164.200 483.800 164.400 ;
        RECT 433.800 163.800 483.800 164.200 ;
        RECT 433.800 163.600 484.200 163.800 ;
        RECT 434.200 163.200 484.200 163.600 ;
        RECT 434.200 163.000 484.600 163.200 ;
        RECT 434.600 162.600 484.600 163.000 ;
        RECT 434.600 162.400 485.000 162.600 ;
        RECT 435.000 162.000 485.000 162.400 ;
        RECT 435.000 161.800 485.400 162.000 ;
        RECT 435.400 161.400 485.400 161.800 ;
        RECT 435.400 161.200 485.800 161.400 ;
        RECT 435.800 160.800 485.800 161.200 ;
        RECT 435.800 160.600 486.200 160.800 ;
        RECT 436.200 160.200 486.200 160.600 ;
        RECT 436.200 160.000 486.600 160.200 ;
        RECT 436.600 159.600 486.600 160.000 ;
        RECT 436.600 159.400 487.000 159.600 ;
        RECT 437.000 159.000 487.000 159.400 ;
        RECT 437.000 158.800 487.400 159.000 ;
        RECT 437.400 158.400 487.400 158.800 ;
        RECT 437.400 158.200 487.800 158.400 ;
        RECT 437.800 157.800 487.800 158.200 ;
        RECT 437.800 157.600 488.200 157.800 ;
        RECT 438.200 157.200 488.200 157.600 ;
        RECT 438.200 157.000 488.600 157.200 ;
        RECT 438.600 156.600 488.600 157.000 ;
        RECT 438.600 156.400 489.000 156.600 ;
        RECT 439.000 156.000 489.000 156.400 ;
        RECT 439.000 155.800 489.400 156.000 ;
        RECT 439.400 155.400 489.400 155.800 ;
        RECT 439.400 155.200 489.800 155.400 ;
        RECT 439.800 154.800 489.800 155.200 ;
        RECT 439.800 154.600 490.200 154.800 ;
        RECT 440.200 154.200 490.200 154.600 ;
        RECT 440.200 154.000 490.600 154.200 ;
        RECT 440.600 153.600 490.600 154.000 ;
        RECT 440.600 153.400 491.000 153.600 ;
        RECT 441.000 153.000 491.000 153.400 ;
        RECT 441.000 152.800 491.400 153.000 ;
        RECT 441.400 152.400 491.400 152.800 ;
        RECT 441.400 152.200 491.800 152.400 ;
        RECT 441.800 151.800 491.800 152.200 ;
        RECT 441.800 151.600 492.200 151.800 ;
        RECT 442.200 151.200 492.200 151.600 ;
        RECT 442.200 151.000 492.600 151.200 ;
        RECT 442.600 150.600 492.600 151.000 ;
        RECT 442.600 150.400 493.000 150.600 ;
        RECT 443.000 150.000 493.000 150.400 ;
        RECT 443.000 149.800 493.400 150.000 ;
        RECT 443.400 149.400 493.400 149.800 ;
        RECT 443.400 149.200 493.800 149.400 ;
        RECT 443.800 148.800 493.800 149.200 ;
        RECT 443.800 148.600 494.200 148.800 ;
        RECT 444.200 148.200 494.200 148.600 ;
        RECT 444.200 148.000 494.600 148.200 ;
        RECT 444.600 147.600 494.600 148.000 ;
        RECT 444.600 147.400 495.000 147.600 ;
        RECT 445.000 147.000 495.000 147.400 ;
        RECT 445.000 146.800 495.400 147.000 ;
        RECT 445.400 146.400 495.400 146.800 ;
        RECT 445.400 146.200 495.800 146.400 ;
        RECT 445.800 145.800 495.800 146.200 ;
        RECT 445.800 145.600 496.200 145.800 ;
        RECT 446.200 145.200 496.200 145.600 ;
        RECT 446.200 145.000 496.600 145.200 ;
        RECT 446.600 144.600 496.600 145.000 ;
        RECT 446.600 144.400 497.000 144.600 ;
        RECT 447.000 144.000 497.000 144.400 ;
        RECT 447.000 143.800 497.400 144.000 ;
        RECT 447.400 143.400 497.400 143.800 ;
        RECT 447.400 143.200 497.800 143.400 ;
        RECT 447.800 142.800 497.800 143.200 ;
        RECT 447.800 142.600 498.200 142.800 ;
        RECT 448.200 142.200 498.200 142.600 ;
        RECT 448.200 142.000 498.600 142.200 ;
        RECT 448.600 141.600 498.600 142.000 ;
        RECT 448.600 141.400 499.000 141.600 ;
        RECT 449.000 141.000 499.000 141.400 ;
        RECT 449.000 140.800 499.400 141.000 ;
        RECT 449.400 140.400 499.400 140.800 ;
        RECT 449.400 140.200 499.800 140.400 ;
        RECT 449.800 139.800 499.800 140.200 ;
        RECT 449.800 139.600 500.200 139.800 ;
        RECT 450.200 139.200 500.200 139.600 ;
        RECT 450.200 139.000 500.600 139.200 ;
        RECT 450.600 138.600 500.600 139.000 ;
        RECT 450.600 138.400 501.000 138.600 ;
        RECT 451.000 138.000 501.000 138.400 ;
        RECT 451.000 137.800 501.400 138.000 ;
        RECT 451.400 137.400 501.400 137.800 ;
        RECT 451.400 137.200 501.800 137.400 ;
        RECT 451.800 136.800 501.800 137.200 ;
        RECT 451.800 136.600 502.200 136.800 ;
        RECT 452.200 136.200 502.200 136.600 ;
        RECT 452.200 136.000 502.600 136.200 ;
        RECT 452.600 135.600 502.600 136.000 ;
        RECT 452.600 135.400 503.000 135.600 ;
        RECT 453.000 135.000 503.000 135.400 ;
        RECT 453.000 134.800 503.400 135.000 ;
        RECT 453.400 134.400 503.400 134.800 ;
        RECT 453.400 134.200 503.800 134.400 ;
        RECT 453.800 133.800 503.800 134.200 ;
        RECT 453.800 133.600 504.200 133.800 ;
        RECT 454.200 133.200 504.200 133.600 ;
        RECT 454.200 133.000 504.600 133.200 ;
        RECT 454.600 132.600 504.600 133.000 ;
        RECT 454.600 132.400 505.000 132.600 ;
        RECT 455.000 132.000 505.000 132.400 ;
        RECT 455.000 131.800 505.400 132.000 ;
        RECT 455.400 131.400 505.400 131.800 ;
        RECT 455.400 131.200 505.800 131.400 ;
        RECT 455.800 130.800 505.800 131.200 ;
        RECT 455.800 130.600 506.200 130.800 ;
        RECT 456.200 130.200 506.200 130.600 ;
        RECT 456.200 130.000 506.600 130.200 ;
        RECT 456.600 129.600 506.600 130.000 ;
        RECT 456.600 129.400 507.000 129.600 ;
        RECT 457.000 129.000 507.000 129.400 ;
        RECT 457.000 128.800 507.400 129.000 ;
        RECT 457.400 128.400 507.400 128.800 ;
        RECT 457.400 128.200 507.800 128.400 ;
        RECT 457.800 127.800 507.800 128.200 ;
        RECT 457.800 127.600 508.200 127.800 ;
        RECT 458.200 127.200 508.200 127.600 ;
        RECT 458.200 127.000 508.600 127.200 ;
        RECT 458.600 126.600 508.600 127.000 ;
        RECT 458.600 126.400 509.000 126.600 ;
        RECT 459.000 126.000 509.000 126.400 ;
        RECT 459.000 125.800 509.400 126.000 ;
        RECT 459.400 125.400 509.400 125.800 ;
        RECT 459.400 125.200 509.800 125.400 ;
        RECT 459.800 124.800 509.800 125.200 ;
        RECT 459.800 124.600 510.200 124.800 ;
        RECT 460.200 124.200 510.200 124.600 ;
        RECT 460.200 124.000 510.600 124.200 ;
        RECT 460.600 123.600 510.600 124.000 ;
        RECT 460.600 123.400 511.000 123.600 ;
        RECT 461.000 123.000 511.000 123.400 ;
        RECT 461.000 122.800 511.400 123.000 ;
        RECT 461.400 122.400 511.400 122.800 ;
        RECT 461.400 122.200 511.800 122.400 ;
        RECT 461.800 121.800 511.800 122.200 ;
        RECT 461.800 121.600 512.200 121.800 ;
        RECT 462.200 121.200 512.200 121.600 ;
        RECT 462.200 121.000 512.600 121.200 ;
        RECT 462.600 120.600 512.600 121.000 ;
        RECT 462.600 120.400 513.000 120.600 ;
        RECT 463.000 120.000 513.000 120.400 ;
        RECT 463.000 119.800 513.400 120.000 ;
        RECT 463.400 119.400 513.400 119.800 ;
        RECT 463.400 119.200 513.800 119.400 ;
        RECT 463.800 118.800 513.800 119.200 ;
        RECT 463.800 118.600 514.200 118.800 ;
        RECT 464.200 118.200 514.200 118.600 ;
        RECT 464.200 118.000 514.600 118.200 ;
        RECT 464.600 117.600 514.600 118.000 ;
        RECT 464.600 117.400 515.000 117.600 ;
        RECT 465.000 117.000 515.000 117.400 ;
        RECT 465.000 116.800 515.400 117.000 ;
        RECT 465.400 116.400 515.400 116.800 ;
        RECT 465.400 116.200 515.800 116.400 ;
        RECT 465.800 115.800 515.800 116.200 ;
        RECT 465.800 115.600 516.200 115.800 ;
        RECT 466.200 115.200 516.200 115.600 ;
        RECT 466.200 115.000 516.600 115.200 ;
        RECT 466.600 114.600 516.600 115.000 ;
        RECT 466.600 114.400 517.000 114.600 ;
        RECT 467.000 114.000 517.000 114.400 ;
        RECT 467.000 113.800 517.400 114.000 ;
        RECT 467.400 113.400 517.400 113.800 ;
        RECT 467.400 113.200 517.800 113.400 ;
        RECT 467.800 112.800 517.800 113.200 ;
        RECT 467.800 112.600 518.200 112.800 ;
        RECT 468.200 112.200 518.200 112.600 ;
        RECT 468.200 112.000 518.600 112.200 ;
        RECT 468.600 111.600 518.600 112.000 ;
        RECT 468.600 111.400 519.000 111.600 ;
        RECT 469.000 111.000 519.000 111.400 ;
        RECT 469.000 110.800 519.400 111.000 ;
        RECT 469.400 110.400 519.400 110.800 ;
        RECT 469.400 110.200 519.800 110.400 ;
        RECT 469.800 109.800 519.800 110.200 ;
        RECT 469.800 109.600 520.200 109.800 ;
        RECT 470.200 109.200 520.200 109.600 ;
        RECT 470.200 109.000 520.600 109.200 ;
        RECT 470.600 108.600 520.600 109.000 ;
        RECT 470.600 108.400 521.000 108.600 ;
        RECT 471.000 108.000 521.000 108.400 ;
        RECT 471.000 107.800 521.400 108.000 ;
        RECT 471.400 107.400 521.400 107.800 ;
        RECT 471.400 107.200 521.800 107.400 ;
        RECT 471.800 106.800 521.800 107.200 ;
        RECT 471.800 106.600 522.200 106.800 ;
        RECT 472.200 106.200 522.200 106.600 ;
        RECT 472.200 106.000 522.600 106.200 ;
        RECT 472.600 105.600 522.600 106.000 ;
        RECT 472.600 105.400 523.000 105.600 ;
        RECT 473.000 105.000 523.000 105.400 ;
        RECT 473.000 104.800 523.400 105.000 ;
        RECT 473.400 104.400 523.400 104.800 ;
        RECT 473.400 104.200 523.800 104.400 ;
        RECT 473.800 103.800 523.800 104.200 ;
        RECT 473.800 103.600 524.200 103.800 ;
        RECT 474.200 103.200 524.200 103.600 ;
        RECT 474.200 103.000 524.600 103.200 ;
        RECT 474.600 102.600 524.600 103.000 ;
        RECT 474.600 102.400 525.000 102.600 ;
        RECT 475.000 102.000 525.000 102.400 ;
        RECT 475.000 101.800 525.400 102.000 ;
        RECT 475.400 101.400 525.400 101.800 ;
        RECT 475.400 101.200 525.800 101.400 ;
        RECT 475.800 100.800 525.800 101.200 ;
        RECT 475.800 100.600 526.200 100.800 ;
        RECT 476.200 100.200 526.200 100.600 ;
        RECT 476.200 100.000 526.600 100.200 ;
        RECT 476.600 99.600 526.600 100.000 ;
        RECT 476.600 99.400 527.000 99.600 ;
        RECT 477.000 99.000 527.000 99.400 ;
        RECT 477.000 98.800 527.400 99.000 ;
        RECT 477.400 98.400 527.400 98.800 ;
        RECT 477.400 98.200 527.800 98.400 ;
        RECT 477.800 97.800 527.800 98.200 ;
        RECT 477.800 97.600 528.200 97.800 ;
        RECT 478.200 97.200 528.200 97.600 ;
        RECT 478.200 97.000 528.600 97.200 ;
        RECT 478.600 96.600 528.600 97.000 ;
        RECT 478.600 96.400 529.000 96.600 ;
        RECT 479.000 96.000 529.000 96.400 ;
        RECT 479.000 95.800 529.400 96.000 ;
        RECT 479.400 95.400 529.400 95.800 ;
        RECT 479.400 95.200 529.800 95.400 ;
        RECT 479.800 94.800 529.800 95.200 ;
        RECT 479.800 94.600 530.200 94.800 ;
        RECT 480.200 94.200 530.200 94.600 ;
        RECT 480.200 94.000 530.600 94.200 ;
        RECT 480.600 93.600 530.600 94.000 ;
        RECT 480.600 93.400 531.000 93.600 ;
        RECT 481.000 93.000 531.000 93.400 ;
        RECT 481.000 92.800 531.400 93.000 ;
        RECT 481.400 92.400 531.400 92.800 ;
        RECT 481.400 92.200 531.800 92.400 ;
        RECT 481.800 91.800 531.800 92.200 ;
        RECT 481.800 91.600 532.200 91.800 ;
        RECT 482.200 91.200 532.200 91.600 ;
        RECT 482.200 91.000 532.600 91.200 ;
        RECT 482.600 90.600 532.600 91.000 ;
        RECT 482.600 90.400 533.000 90.600 ;
        RECT 483.000 90.000 533.000 90.400 ;
        RECT 483.000 89.800 533.400 90.000 ;
        RECT 483.400 89.400 533.400 89.800 ;
        RECT 483.400 89.200 533.800 89.400 ;
        RECT 483.800 88.800 533.800 89.200 ;
        RECT 483.800 88.600 534.200 88.800 ;
        RECT 484.200 88.200 534.200 88.600 ;
        RECT 484.200 88.000 534.600 88.200 ;
        RECT 484.600 87.600 534.600 88.000 ;
        RECT 535.000 87.600 585.000 342.600 ;
        RECT 484.600 87.400 585.000 87.600 ;
        RECT 485.000 86.800 585.000 87.400 ;
        RECT 485.400 86.200 585.000 86.800 ;
        RECT 485.800 85.600 585.000 86.200 ;
        RECT 486.200 85.000 585.000 85.600 ;
        RECT 486.600 84.400 585.000 85.000 ;
        RECT 487.000 83.800 585.000 84.400 ;
        RECT 487.400 83.200 585.000 83.800 ;
        RECT 487.800 82.600 585.000 83.200 ;
        RECT 488.200 82.000 585.000 82.600 ;
        RECT 488.600 81.400 585.000 82.000 ;
        RECT 489.000 80.800 585.000 81.400 ;
        RECT 489.400 80.200 585.000 80.800 ;
        RECT 489.800 79.600 585.000 80.200 ;
        RECT 490.200 79.000 585.000 79.600 ;
        RECT 490.600 78.400 585.000 79.000 ;
        RECT 491.000 77.800 585.000 78.400 ;
        RECT 491.400 77.200 585.000 77.800 ;
        RECT 491.800 76.600 585.000 77.200 ;
        RECT 492.200 76.000 585.000 76.600 ;
        RECT 492.600 75.400 585.000 76.000 ;
        RECT 493.000 74.800 585.000 75.400 ;
        RECT 493.400 74.200 585.000 74.800 ;
        RECT 493.800 73.600 585.000 74.200 ;
        RECT 494.200 73.000 585.000 73.600 ;
        RECT 494.600 72.400 585.000 73.000 ;
        RECT 495.000 71.800 585.000 72.400 ;
        RECT 495.400 71.200 585.000 71.800 ;
        RECT 495.800 70.600 585.000 71.200 ;
        RECT 496.200 70.000 585.000 70.600 ;
        RECT 496.600 69.400 585.000 70.000 ;
        RECT 497.000 68.800 585.000 69.400 ;
        RECT 497.400 68.200 585.000 68.800 ;
        RECT 497.800 67.600 585.000 68.200 ;
        RECT 498.200 67.000 585.000 67.600 ;
        RECT 498.600 66.400 585.000 67.000 ;
        RECT 499.000 65.800 585.000 66.400 ;
        RECT 499.400 65.200 585.000 65.800 ;
        RECT 499.800 64.600 585.000 65.200 ;
        RECT 500.200 64.000 585.000 64.600 ;
        RECT 500.600 63.400 585.000 64.000 ;
        RECT 501.000 62.800 585.000 63.400 ;
        RECT 501.400 62.200 585.000 62.800 ;
        RECT 501.800 61.600 585.000 62.200 ;
        RECT 502.200 61.000 585.000 61.600 ;
        RECT 502.600 60.400 585.000 61.000 ;
        RECT 503.000 59.800 585.000 60.400 ;
        RECT 503.400 59.200 585.000 59.800 ;
        RECT 503.800 58.600 585.000 59.200 ;
        RECT 504.200 58.000 585.000 58.600 ;
        RECT 504.600 57.400 585.000 58.000 ;
        RECT 505.000 56.800 585.000 57.400 ;
        RECT 505.400 56.200 585.000 56.800 ;
        RECT 505.800 55.600 585.000 56.200 ;
        RECT 506.200 55.000 585.000 55.600 ;
        RECT 506.600 54.400 585.000 55.000 ;
        RECT 507.000 53.800 585.000 54.400 ;
        RECT 507.400 53.200 585.000 53.800 ;
        RECT 507.800 52.600 585.000 53.200 ;
        RECT 508.200 52.000 585.000 52.600 ;
        RECT 508.600 51.400 585.000 52.000 ;
        RECT 509.000 50.800 585.000 51.400 ;
        RECT 509.400 50.200 585.000 50.800 ;
        RECT 509.800 49.600 585.000 50.200 ;
        RECT 510.200 49.000 585.000 49.600 ;
        RECT 510.600 48.400 585.000 49.000 ;
        RECT 511.000 47.800 585.000 48.400 ;
        RECT 511.400 47.200 585.000 47.800 ;
        RECT 511.800 46.600 585.000 47.200 ;
        RECT 512.200 46.000 585.000 46.600 ;
        RECT 512.600 45.400 585.000 46.000 ;
        RECT 513.000 44.800 585.000 45.400 ;
        RECT 513.400 44.200 585.000 44.800 ;
        RECT 513.800 43.600 585.000 44.200 ;
        RECT 514.200 43.000 585.000 43.600 ;
        RECT 514.600 42.400 585.000 43.000 ;
        RECT 515.000 41.800 585.000 42.400 ;
        RECT 515.400 41.200 585.000 41.800 ;
        RECT 515.800 40.600 585.000 41.200 ;
        RECT 516.200 40.000 585.000 40.600 ;
        RECT 516.600 39.400 585.000 40.000 ;
        RECT 517.000 38.800 585.000 39.400 ;
        RECT 517.400 38.200 585.000 38.800 ;
        RECT 517.800 37.600 585.000 38.200 ;
        RECT 518.200 37.000 585.000 37.600 ;
        RECT 518.600 36.400 585.000 37.000 ;
        RECT 519.000 35.800 585.000 36.400 ;
        RECT 519.400 35.200 585.000 35.800 ;
        RECT 519.800 34.600 585.000 35.200 ;
        RECT 520.200 34.000 585.000 34.600 ;
        RECT 520.600 33.400 585.000 34.000 ;
        RECT 521.000 32.800 585.000 33.400 ;
        RECT 521.400 32.200 585.000 32.800 ;
        RECT 521.800 31.600 585.000 32.200 ;
        RECT 522.200 31.000 585.000 31.600 ;
        RECT 522.600 30.400 585.000 31.000 ;
        RECT 523.000 29.800 585.000 30.400 ;
        RECT 523.400 29.200 585.000 29.800 ;
        RECT 523.800 28.600 585.000 29.200 ;
        RECT 524.200 28.000 585.000 28.600 ;
        RECT 524.600 27.400 585.000 28.000 ;
        RECT 525.000 26.800 585.000 27.400 ;
        RECT 525.400 26.200 585.000 26.800 ;
        RECT 525.800 25.600 585.000 26.200 ;
        RECT 526.200 25.000 585.000 25.600 ;
        RECT 526.600 24.400 585.000 25.000 ;
        RECT 527.000 23.800 585.000 24.400 ;
        RECT 527.400 23.200 585.000 23.800 ;
        RECT 527.800 22.600 585.000 23.200 ;
        RECT 528.200 22.000 585.000 22.600 ;
        RECT 528.600 21.400 585.000 22.000 ;
        RECT 529.000 20.800 585.000 21.400 ;
        RECT 529.400 20.200 585.000 20.800 ;
        RECT 529.800 19.600 585.000 20.200 ;
        RECT 530.200 19.000 585.000 19.600 ;
        RECT 530.600 18.400 585.000 19.000 ;
        RECT 531.000 17.800 585.000 18.400 ;
        RECT 531.400 17.200 585.000 17.800 ;
        RECT 531.800 16.600 585.000 17.200 ;
        RECT 532.200 16.000 585.000 16.600 ;
        RECT 532.600 15.400 585.000 16.000 ;
        RECT 533.000 14.800 585.000 15.400 ;
        RECT 533.400 14.200 585.000 14.800 ;
        RECT 533.800 13.600 585.000 14.200 ;
        RECT 534.200 13.000 585.000 13.600 ;
        RECT 534.600 12.400 585.000 13.000 ;
    END
  END vss
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 1200.000 352.200 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 1200.000 352.200 ;
      LAYER Metal4 ;
        RECT 0.000 0.000 1200.000 352.200 ;
      LAYER Metal5 ;
        RECT 725.000 342.000 775.000 342.600 ;
        RECT 915.000 342.000 965.000 342.600 ;
        RECT 724.800 341.400 775.200 342.000 ;
        RECT 915.000 341.400 965.400 342.000 ;
        RECT 724.600 340.800 775.400 341.400 ;
        RECT 915.000 340.800 965.800 341.400 ;
        RECT 724.300 340.200 775.700 340.800 ;
        RECT 915.000 340.200 966.200 340.800 ;
        RECT 724.100 339.600 775.900 340.200 ;
        RECT 915.000 339.600 966.600 340.200 ;
        RECT 723.900 339.000 776.100 339.600 ;
        RECT 915.000 339.000 967.000 339.600 ;
        RECT 723.600 338.400 776.400 339.000 ;
        RECT 915.000 338.400 967.400 339.000 ;
        RECT 723.400 337.800 776.600 338.400 ;
        RECT 915.000 337.800 967.800 338.400 ;
        RECT 723.200 337.200 776.800 337.800 ;
        RECT 915.000 337.200 968.200 337.800 ;
        RECT 723.000 336.600 777.000 337.200 ;
        RECT 915.000 336.600 968.600 337.200 ;
        RECT 722.800 336.000 777.200 336.600 ;
        RECT 915.000 336.000 969.000 336.600 ;
        RECT 722.500 335.400 777.500 336.000 ;
        RECT 915.000 335.400 969.400 336.000 ;
        RECT 722.300 334.800 777.700 335.400 ;
        RECT 915.000 334.800 969.800 335.400 ;
        RECT 722.100 334.200 777.900 334.800 ;
        RECT 915.000 334.200 970.200 334.800 ;
        RECT 721.800 333.600 778.200 334.200 ;
        RECT 915.000 333.600 970.600 334.200 ;
        RECT 721.600 333.000 778.400 333.600 ;
        RECT 915.000 333.000 971.000 333.600 ;
        RECT 721.400 332.400 778.600 333.000 ;
        RECT 915.000 332.400 971.400 333.000 ;
        RECT 721.200 331.800 778.800 332.400 ;
        RECT 915.000 331.800 971.800 332.400 ;
        RECT 721.000 331.200 779.000 331.800 ;
        RECT 915.000 331.200 972.200 331.800 ;
        RECT 720.700 330.600 779.300 331.200 ;
        RECT 915.000 330.600 972.600 331.200 ;
        RECT 720.500 330.000 779.500 330.600 ;
        RECT 915.000 330.000 973.000 330.600 ;
        RECT 720.300 329.400 779.700 330.000 ;
        RECT 915.000 329.400 973.400 330.000 ;
        RECT 720.000 328.800 780.000 329.400 ;
        RECT 915.000 328.800 973.800 329.400 ;
        RECT 719.800 328.200 780.200 328.800 ;
        RECT 915.000 328.200 974.200 328.800 ;
        RECT 719.600 327.600 780.400 328.200 ;
        RECT 915.000 327.600 974.600 328.200 ;
        RECT 719.400 327.000 780.600 327.600 ;
        RECT 915.000 327.000 975.000 327.600 ;
        RECT 719.200 326.400 780.800 327.000 ;
        RECT 915.000 326.400 975.400 327.000 ;
        RECT 718.900 325.800 781.100 326.400 ;
        RECT 915.000 325.800 975.800 326.400 ;
        RECT 718.700 325.200 781.300 325.800 ;
        RECT 915.000 325.200 976.200 325.800 ;
        RECT 718.500 324.600 781.500 325.200 ;
        RECT 915.000 324.600 976.600 325.200 ;
        RECT 718.200 324.000 781.800 324.600 ;
        RECT 915.000 324.000 977.000 324.600 ;
        RECT 718.000 323.400 782.000 324.000 ;
        RECT 915.000 323.400 977.400 324.000 ;
        RECT 717.800 322.800 782.200 323.400 ;
        RECT 915.000 322.800 977.800 323.400 ;
        RECT 717.600 322.200 782.400 322.800 ;
        RECT 915.000 322.200 978.200 322.800 ;
        RECT 717.400 321.600 782.600 322.200 ;
        RECT 915.000 321.600 978.600 322.200 ;
        RECT 717.100 321.000 782.900 321.600 ;
        RECT 915.000 321.000 979.000 321.600 ;
        RECT 716.900 320.400 783.100 321.000 ;
        RECT 915.000 320.400 979.400 321.000 ;
        RECT 716.700 319.800 783.300 320.400 ;
        RECT 915.000 319.800 979.800 320.400 ;
        RECT 716.400 319.200 783.600 319.800 ;
        RECT 915.000 319.200 980.200 319.800 ;
        RECT 716.200 318.600 783.800 319.200 ;
        RECT 915.000 318.600 980.600 319.200 ;
        RECT 716.000 318.000 784.000 318.600 ;
        RECT 915.000 318.000 981.000 318.600 ;
        RECT 715.800 317.400 784.200 318.000 ;
        RECT 915.000 317.400 981.400 318.000 ;
        RECT 715.600 316.800 784.400 317.400 ;
        RECT 915.000 316.800 981.800 317.400 ;
        RECT 715.300 316.200 784.700 316.800 ;
        RECT 915.000 316.200 982.200 316.800 ;
        RECT 715.100 315.600 784.900 316.200 ;
        RECT 915.000 315.600 982.600 316.200 ;
        RECT 714.900 315.000 785.100 315.600 ;
        RECT 915.000 315.000 983.000 315.600 ;
        RECT 714.600 314.400 785.400 315.000 ;
        RECT 915.000 314.400 983.400 315.000 ;
        RECT 714.400 313.800 785.600 314.400 ;
        RECT 915.000 313.800 983.800 314.400 ;
        RECT 714.200 313.200 785.800 313.800 ;
        RECT 915.000 313.200 984.200 313.800 ;
        RECT 714.000 312.600 786.000 313.200 ;
        RECT 915.000 312.600 984.600 313.200 ;
        RECT 713.800 312.000 786.200 312.600 ;
        RECT 915.000 312.000 985.000 312.600 ;
        RECT 713.500 311.400 786.500 312.000 ;
        RECT 915.000 311.400 985.400 312.000 ;
        RECT 713.300 310.800 786.700 311.400 ;
        RECT 915.000 310.800 985.800 311.400 ;
        RECT 713.100 310.200 786.900 310.800 ;
        RECT 915.000 310.200 986.200 310.800 ;
        RECT 712.800 309.600 787.200 310.200 ;
        RECT 915.000 309.600 986.600 310.200 ;
        RECT 712.600 309.000 787.400 309.600 ;
        RECT 915.000 309.000 987.000 309.600 ;
        RECT 712.400 308.400 787.600 309.000 ;
        RECT 915.000 308.400 987.400 309.000 ;
        RECT 712.200 307.800 787.800 308.400 ;
        RECT 915.000 307.800 987.800 308.400 ;
        RECT 712.000 307.200 788.000 307.800 ;
        RECT 915.000 307.200 988.200 307.800 ;
        RECT 711.700 306.600 788.300 307.200 ;
        RECT 915.000 306.600 988.600 307.200 ;
        RECT 711.500 306.000 788.500 306.600 ;
        RECT 915.000 306.000 989.000 306.600 ;
        RECT 711.300 305.400 788.700 306.000 ;
        RECT 915.000 305.400 989.400 306.000 ;
        RECT 711.000 304.800 789.000 305.400 ;
        RECT 915.000 304.800 989.800 305.400 ;
        RECT 710.800 304.200 789.200 304.800 ;
        RECT 915.000 304.200 990.200 304.800 ;
        RECT 710.600 303.600 789.400 304.200 ;
        RECT 915.000 303.600 990.600 304.200 ;
        RECT 710.400 303.000 789.600 303.600 ;
        RECT 915.000 303.000 991.000 303.600 ;
        RECT 710.200 302.400 789.800 303.000 ;
        RECT 915.000 302.400 991.400 303.000 ;
        RECT 709.900 301.800 790.100 302.400 ;
        RECT 915.000 301.800 991.800 302.400 ;
        RECT 709.700 301.200 790.300 301.800 ;
        RECT 915.000 301.200 992.200 301.800 ;
        RECT 709.500 300.600 790.500 301.200 ;
        RECT 915.000 300.600 992.600 301.200 ;
        RECT 709.200 300.000 790.800 300.600 ;
        RECT 915.000 300.000 993.000 300.600 ;
        RECT 709.000 299.400 791.000 300.000 ;
        RECT 915.000 299.400 993.400 300.000 ;
        RECT 708.800 298.800 791.200 299.400 ;
        RECT 915.000 298.800 993.800 299.400 ;
        RECT 708.600 298.200 791.400 298.800 ;
        RECT 915.000 298.200 994.200 298.800 ;
        RECT 708.400 297.600 791.600 298.200 ;
        RECT 915.000 297.600 994.600 298.200 ;
        RECT 708.100 297.000 791.900 297.600 ;
        RECT 915.000 297.000 995.000 297.600 ;
        RECT 707.900 296.400 792.100 297.000 ;
        RECT 915.000 296.400 995.400 297.000 ;
        RECT 707.700 295.800 792.300 296.400 ;
        RECT 915.000 295.800 995.800 296.400 ;
        RECT 707.400 295.200 792.600 295.800 ;
        RECT 915.000 295.200 996.200 295.800 ;
        RECT 707.200 294.600 792.800 295.200 ;
        RECT 915.000 294.600 996.600 295.200 ;
        RECT 707.000 294.000 793.000 294.600 ;
        RECT 915.000 294.000 997.000 294.600 ;
        RECT 706.800 293.400 793.200 294.000 ;
        RECT 915.000 293.400 997.400 294.000 ;
        RECT 706.600 292.800 793.400 293.400 ;
        RECT 915.000 292.800 997.800 293.400 ;
        RECT 706.300 292.200 793.700 292.800 ;
        RECT 915.000 292.200 998.200 292.800 ;
        RECT 706.100 291.600 793.900 292.200 ;
        RECT 915.000 291.600 998.600 292.200 ;
        RECT 705.900 291.000 794.100 291.600 ;
        RECT 915.000 291.000 999.000 291.600 ;
        RECT 705.600 290.400 794.400 291.000 ;
        RECT 915.000 290.400 999.400 291.000 ;
        RECT 705.400 289.800 794.600 290.400 ;
        RECT 915.000 289.800 999.800 290.400 ;
        RECT 705.200 289.200 794.800 289.800 ;
        RECT 915.000 289.200 1000.200 289.800 ;
        RECT 705.000 288.600 795.000 289.200 ;
        RECT 915.000 288.600 1000.600 289.200 ;
        RECT 704.800 288.000 795.200 288.600 ;
        RECT 915.000 288.000 1001.000 288.600 ;
        RECT 704.500 287.400 795.500 288.000 ;
        RECT 915.000 287.400 1001.400 288.000 ;
        RECT 704.300 286.800 795.700 287.400 ;
        RECT 915.000 286.800 1001.800 287.400 ;
        RECT 704.100 286.200 795.900 286.800 ;
        RECT 915.000 286.200 1002.200 286.800 ;
        RECT 703.800 285.600 796.200 286.200 ;
        RECT 915.000 285.600 1002.600 286.200 ;
        RECT 703.600 285.000 796.400 285.600 ;
        RECT 915.000 285.000 1003.000 285.600 ;
        RECT 703.400 284.400 796.600 285.000 ;
        RECT 915.000 284.400 1003.400 285.000 ;
        RECT 703.200 283.800 796.800 284.400 ;
        RECT 915.000 283.800 1003.800 284.400 ;
        RECT 703.000 283.200 797.000 283.800 ;
        RECT 915.000 283.200 1004.200 283.800 ;
        RECT 702.700 282.600 797.300 283.200 ;
        RECT 915.000 282.600 1004.600 283.200 ;
        RECT 702.500 282.000 797.500 282.600 ;
        RECT 915.000 282.000 1005.000 282.600 ;
        RECT 702.300 281.400 797.700 282.000 ;
        RECT 915.000 281.400 1005.400 282.000 ;
        RECT 702.000 280.800 798.000 281.400 ;
        RECT 915.000 280.800 1005.800 281.400 ;
        RECT 701.800 280.200 798.200 280.800 ;
        RECT 915.000 280.200 1006.200 280.800 ;
        RECT 701.600 279.600 798.400 280.200 ;
        RECT 915.000 279.600 1006.600 280.200 ;
        RECT 701.400 279.000 798.600 279.600 ;
        RECT 915.000 279.000 1007.000 279.600 ;
        RECT 701.200 278.400 798.800 279.000 ;
        RECT 915.000 278.400 1007.400 279.000 ;
        RECT 700.900 277.800 799.100 278.400 ;
        RECT 915.000 277.800 1007.800 278.400 ;
        RECT 700.700 277.200 799.300 277.800 ;
        RECT 915.000 277.200 1008.200 277.800 ;
        RECT 700.500 276.600 799.500 277.200 ;
        RECT 915.000 276.600 1008.600 277.200 ;
        RECT 700.200 276.000 799.800 276.600 ;
        RECT 915.000 276.000 1009.000 276.600 ;
        RECT 700.000 275.400 800.000 276.000 ;
        RECT 915.000 275.400 1009.400 276.000 ;
        RECT 699.800 275.200 800.200 275.400 ;
        RECT 699.800 274.800 749.800 275.200 ;
        RECT 699.600 274.600 749.800 274.800 ;
        RECT 750.200 274.800 800.200 275.200 ;
        RECT 915.000 274.800 1009.800 275.400 ;
        RECT 750.200 274.600 800.400 274.800 ;
        RECT 699.600 274.200 749.600 274.600 ;
        RECT 699.400 274.000 749.600 274.200 ;
        RECT 750.400 274.200 800.400 274.600 ;
        RECT 915.000 274.200 1010.200 274.800 ;
        RECT 750.400 274.000 800.600 274.200 ;
        RECT 699.400 273.600 749.400 274.000 ;
        RECT 699.100 273.400 749.400 273.600 ;
        RECT 750.600 273.600 800.600 274.000 ;
        RECT 915.000 273.600 1010.600 274.200 ;
        RECT 750.600 273.400 800.900 273.600 ;
        RECT 699.100 273.000 749.100 273.400 ;
        RECT 698.900 272.800 749.100 273.000 ;
        RECT 750.900 273.000 800.900 273.400 ;
        RECT 915.000 273.000 1011.000 273.600 ;
        RECT 750.900 272.800 801.100 273.000 ;
        RECT 698.900 272.400 748.900 272.800 ;
        RECT 698.700 272.200 748.900 272.400 ;
        RECT 751.100 272.400 801.100 272.800 ;
        RECT 915.000 272.400 1011.400 273.000 ;
        RECT 751.100 272.200 801.300 272.400 ;
        RECT 698.700 271.800 748.700 272.200 ;
        RECT 698.400 271.600 748.700 271.800 ;
        RECT 751.300 271.800 801.300 272.200 ;
        RECT 915.000 271.800 1011.800 272.400 ;
        RECT 751.300 271.600 801.600 271.800 ;
        RECT 698.400 271.200 748.400 271.600 ;
        RECT 698.200 271.000 748.400 271.200 ;
        RECT 751.600 271.200 801.600 271.600 ;
        RECT 915.000 271.200 1012.200 271.800 ;
        RECT 751.600 271.000 801.800 271.200 ;
        RECT 698.200 270.600 748.200 271.000 ;
        RECT 698.000 270.400 748.200 270.600 ;
        RECT 751.800 270.600 801.800 271.000 ;
        RECT 915.000 270.600 1012.600 271.200 ;
        RECT 751.800 270.400 802.000 270.600 ;
        RECT 698.000 270.000 748.000 270.400 ;
        RECT 697.800 269.800 748.000 270.000 ;
        RECT 752.000 270.000 802.000 270.400 ;
        RECT 915.000 270.000 1013.000 270.600 ;
        RECT 752.000 269.800 802.200 270.000 ;
        RECT 697.800 269.400 747.800 269.800 ;
        RECT 697.600 269.200 747.800 269.400 ;
        RECT 752.200 269.400 802.200 269.800 ;
        RECT 915.000 269.400 1013.400 270.000 ;
        RECT 752.200 269.200 802.400 269.400 ;
        RECT 697.600 268.800 747.600 269.200 ;
        RECT 697.300 268.600 747.600 268.800 ;
        RECT 752.400 268.800 802.400 269.200 ;
        RECT 915.000 268.800 1013.800 269.400 ;
        RECT 752.400 268.600 802.700 268.800 ;
        RECT 697.300 268.200 747.300 268.600 ;
        RECT 697.100 268.000 747.300 268.200 ;
        RECT 752.700 268.200 802.700 268.600 ;
        RECT 915.000 268.200 1014.200 268.800 ;
        RECT 752.700 268.000 802.900 268.200 ;
        RECT 697.100 267.600 747.100 268.000 ;
        RECT 696.900 267.400 747.100 267.600 ;
        RECT 752.900 267.600 802.900 268.000 ;
        RECT 915.000 267.600 1014.600 268.200 ;
        RECT 752.900 267.400 803.100 267.600 ;
        RECT 696.900 267.000 746.900 267.400 ;
        RECT 696.600 266.800 746.900 267.000 ;
        RECT 753.100 267.000 803.100 267.400 ;
        RECT 915.000 267.000 1015.000 267.600 ;
        RECT 753.100 266.800 803.400 267.000 ;
        RECT 696.600 266.400 746.600 266.800 ;
        RECT 696.400 266.200 746.600 266.400 ;
        RECT 753.400 266.400 803.400 266.800 ;
        RECT 915.000 266.800 1015.400 267.000 ;
        RECT 753.400 266.200 803.600 266.400 ;
        RECT 696.400 265.800 746.400 266.200 ;
        RECT 696.200 265.600 746.400 265.800 ;
        RECT 753.600 265.800 803.600 266.200 ;
        RECT 753.600 265.600 803.800 265.800 ;
        RECT 696.200 265.200 746.200 265.600 ;
        RECT 696.000 265.000 746.200 265.200 ;
        RECT 753.800 265.200 803.800 265.600 ;
        RECT 753.800 265.000 804.000 265.200 ;
        RECT 696.000 264.600 746.000 265.000 ;
        RECT 695.800 264.400 746.000 264.600 ;
        RECT 754.000 264.600 804.000 265.000 ;
        RECT 754.000 264.400 804.200 264.600 ;
        RECT 695.800 264.000 745.800 264.400 ;
        RECT 695.500 263.800 745.800 264.000 ;
        RECT 754.200 264.000 804.200 264.400 ;
        RECT 754.200 263.800 804.500 264.000 ;
        RECT 695.500 263.400 745.500 263.800 ;
        RECT 695.300 263.200 745.500 263.400 ;
        RECT 754.500 263.400 804.500 263.800 ;
        RECT 754.500 263.200 804.700 263.400 ;
        RECT 695.300 262.800 745.300 263.200 ;
        RECT 695.100 262.600 745.300 262.800 ;
        RECT 754.700 262.800 804.700 263.200 ;
        RECT 754.700 262.600 804.900 262.800 ;
        RECT 695.100 262.200 745.100 262.600 ;
        RECT 694.800 262.000 745.100 262.200 ;
        RECT 754.900 262.200 804.900 262.600 ;
        RECT 754.900 262.000 805.200 262.200 ;
        RECT 694.800 261.600 744.800 262.000 ;
        RECT 694.600 261.400 744.800 261.600 ;
        RECT 755.200 261.600 805.200 262.000 ;
        RECT 755.200 261.400 805.400 261.600 ;
        RECT 694.600 261.000 744.600 261.400 ;
        RECT 694.400 260.800 744.600 261.000 ;
        RECT 755.400 261.000 805.400 261.400 ;
        RECT 755.400 260.800 805.600 261.000 ;
        RECT 694.400 260.400 744.400 260.800 ;
        RECT 694.200 260.200 744.400 260.400 ;
        RECT 755.600 260.400 805.600 260.800 ;
        RECT 755.600 260.200 805.800 260.400 ;
        RECT 694.200 259.800 744.200 260.200 ;
        RECT 694.000 259.600 744.200 259.800 ;
        RECT 755.800 259.800 805.800 260.200 ;
        RECT 755.800 259.600 806.000 259.800 ;
        RECT 694.000 259.200 744.000 259.600 ;
        RECT 693.700 259.000 744.000 259.200 ;
        RECT 756.000 259.200 806.000 259.600 ;
        RECT 756.000 259.000 806.300 259.200 ;
        RECT 693.700 258.600 743.700 259.000 ;
        RECT 693.500 258.400 743.700 258.600 ;
        RECT 756.300 258.600 806.300 259.000 ;
        RECT 756.300 258.400 806.500 258.600 ;
        RECT 693.500 258.000 743.500 258.400 ;
        RECT 693.300 257.800 743.500 258.000 ;
        RECT 756.500 258.000 806.500 258.400 ;
        RECT 756.500 257.800 806.700 258.000 ;
        RECT 693.300 257.400 743.300 257.800 ;
        RECT 693.000 257.200 743.300 257.400 ;
        RECT 756.700 257.400 806.700 257.800 ;
        RECT 756.700 257.200 807.000 257.400 ;
        RECT 693.000 256.800 743.000 257.200 ;
        RECT 692.800 256.600 743.000 256.800 ;
        RECT 757.000 256.800 807.000 257.200 ;
        RECT 757.000 256.600 807.200 256.800 ;
        RECT 692.800 256.200 742.800 256.600 ;
        RECT 692.600 256.000 742.800 256.200 ;
        RECT 757.200 256.200 807.200 256.600 ;
        RECT 757.200 256.000 807.400 256.200 ;
        RECT 692.600 255.600 742.600 256.000 ;
        RECT 692.400 255.400 742.600 255.600 ;
        RECT 757.400 255.600 807.400 256.000 ;
        RECT 757.400 255.400 807.600 255.600 ;
        RECT 692.400 255.000 742.400 255.400 ;
        RECT 692.200 254.800 742.400 255.000 ;
        RECT 757.600 255.000 807.600 255.400 ;
        RECT 757.600 254.800 807.800 255.000 ;
        RECT 692.200 254.400 742.200 254.800 ;
        RECT 691.900 254.200 742.200 254.400 ;
        RECT 757.800 254.400 807.800 254.800 ;
        RECT 757.800 254.200 808.100 254.400 ;
        RECT 691.900 253.800 741.900 254.200 ;
        RECT 691.700 253.600 741.900 253.800 ;
        RECT 758.100 253.800 808.100 254.200 ;
        RECT 758.100 253.600 808.300 253.800 ;
        RECT 691.700 253.200 741.700 253.600 ;
        RECT 691.500 253.000 741.700 253.200 ;
        RECT 758.300 253.200 808.300 253.600 ;
        RECT 758.300 253.000 808.500 253.200 ;
        RECT 691.500 252.600 741.500 253.000 ;
        RECT 691.200 252.400 741.500 252.600 ;
        RECT 758.500 252.600 808.500 253.000 ;
        RECT 758.500 252.400 808.800 252.600 ;
        RECT 691.200 252.000 741.200 252.400 ;
        RECT 691.000 251.800 741.200 252.000 ;
        RECT 758.800 252.000 808.800 252.400 ;
        RECT 758.800 251.800 809.000 252.000 ;
        RECT 691.000 251.400 741.000 251.800 ;
        RECT 690.800 251.200 741.000 251.400 ;
        RECT 759.000 251.400 809.000 251.800 ;
        RECT 759.000 251.200 809.200 251.400 ;
        RECT 690.800 250.800 740.800 251.200 ;
        RECT 690.600 250.600 740.800 250.800 ;
        RECT 759.200 250.800 809.200 251.200 ;
        RECT 759.200 250.600 809.400 250.800 ;
        RECT 690.600 250.200 740.600 250.600 ;
        RECT 690.400 250.000 740.600 250.200 ;
        RECT 759.400 250.200 809.400 250.600 ;
        RECT 759.400 250.000 809.600 250.200 ;
        RECT 690.400 249.600 740.400 250.000 ;
        RECT 690.100 249.400 740.400 249.600 ;
        RECT 759.600 249.600 809.600 250.000 ;
        RECT 759.600 249.400 809.900 249.600 ;
        RECT 690.100 249.000 740.100 249.400 ;
        RECT 689.900 248.800 740.100 249.000 ;
        RECT 759.900 249.000 809.900 249.400 ;
        RECT 759.900 248.800 810.100 249.000 ;
        RECT 689.900 248.400 739.900 248.800 ;
        RECT 689.700 248.200 739.900 248.400 ;
        RECT 760.100 248.400 810.100 248.800 ;
        RECT 760.100 248.200 810.300 248.400 ;
        RECT 689.700 247.800 739.700 248.200 ;
        RECT 689.400 247.600 739.700 247.800 ;
        RECT 760.300 247.800 810.300 248.200 ;
        RECT 760.300 247.600 810.600 247.800 ;
        RECT 689.400 247.200 739.400 247.600 ;
        RECT 689.200 247.000 739.400 247.200 ;
        RECT 760.600 247.200 810.600 247.600 ;
        RECT 760.600 247.000 810.800 247.200 ;
        RECT 689.200 246.600 739.200 247.000 ;
        RECT 689.000 246.400 739.200 246.600 ;
        RECT 760.800 246.600 810.800 247.000 ;
        RECT 760.800 246.400 811.000 246.600 ;
        RECT 689.000 246.000 739.000 246.400 ;
        RECT 688.800 245.800 739.000 246.000 ;
        RECT 761.000 246.000 811.000 246.400 ;
        RECT 761.000 245.800 811.200 246.000 ;
        RECT 688.800 245.400 738.800 245.800 ;
        RECT 688.600 245.200 738.800 245.400 ;
        RECT 761.200 245.400 811.200 245.800 ;
        RECT 761.200 245.200 811.400 245.400 ;
        RECT 688.600 244.800 738.600 245.200 ;
        RECT 688.300 244.600 738.600 244.800 ;
        RECT 761.400 244.800 811.400 245.200 ;
        RECT 761.400 244.600 811.700 244.800 ;
        RECT 688.300 244.200 738.300 244.600 ;
        RECT 688.100 244.000 738.300 244.200 ;
        RECT 761.700 244.200 811.700 244.600 ;
        RECT 761.700 244.000 811.900 244.200 ;
        RECT 688.100 243.600 738.100 244.000 ;
        RECT 687.900 243.400 738.100 243.600 ;
        RECT 761.900 243.600 811.900 244.000 ;
        RECT 761.900 243.400 812.100 243.600 ;
        RECT 687.900 243.000 737.900 243.400 ;
        RECT 687.600 242.800 737.900 243.000 ;
        RECT 762.100 243.000 812.100 243.400 ;
        RECT 762.100 242.800 812.400 243.000 ;
        RECT 687.600 242.400 737.600 242.800 ;
        RECT 687.400 242.200 737.600 242.400 ;
        RECT 762.400 242.400 812.400 242.800 ;
        RECT 762.400 242.200 812.600 242.400 ;
        RECT 687.400 241.800 737.400 242.200 ;
        RECT 687.200 241.600 737.400 241.800 ;
        RECT 762.600 241.800 812.600 242.200 ;
        RECT 762.600 241.600 812.800 241.800 ;
        RECT 687.200 241.200 737.200 241.600 ;
        RECT 687.000 241.000 737.200 241.200 ;
        RECT 762.800 241.200 812.800 241.600 ;
        RECT 762.800 241.000 813.000 241.200 ;
        RECT 687.000 240.600 737.000 241.000 ;
        RECT 686.800 240.400 737.000 240.600 ;
        RECT 763.000 240.600 813.000 241.000 ;
        RECT 763.000 240.400 813.200 240.600 ;
        RECT 686.800 240.000 736.800 240.400 ;
        RECT 686.500 239.800 736.800 240.000 ;
        RECT 763.200 240.000 813.200 240.400 ;
        RECT 763.200 239.800 813.500 240.000 ;
        RECT 686.500 239.400 736.500 239.800 ;
        RECT 686.300 239.200 736.500 239.400 ;
        RECT 763.500 239.400 813.500 239.800 ;
        RECT 763.500 239.200 813.700 239.400 ;
        RECT 686.300 238.800 736.300 239.200 ;
        RECT 686.100 238.600 736.300 238.800 ;
        RECT 763.700 238.800 813.700 239.200 ;
        RECT 763.700 238.600 813.900 238.800 ;
        RECT 686.100 238.200 736.100 238.600 ;
        RECT 685.800 238.000 736.100 238.200 ;
        RECT 763.900 238.200 813.900 238.600 ;
        RECT 763.900 238.000 814.200 238.200 ;
        RECT 685.800 237.600 735.800 238.000 ;
        RECT 685.600 237.400 735.800 237.600 ;
        RECT 764.200 237.600 814.200 238.000 ;
        RECT 764.200 237.400 814.400 237.600 ;
        RECT 685.600 237.000 735.600 237.400 ;
        RECT 685.400 236.800 735.600 237.000 ;
        RECT 764.400 237.000 814.400 237.400 ;
        RECT 764.400 236.800 814.600 237.000 ;
        RECT 685.400 236.400 735.400 236.800 ;
        RECT 685.200 236.200 735.400 236.400 ;
        RECT 764.600 236.400 814.600 236.800 ;
        RECT 764.600 236.200 814.800 236.400 ;
        RECT 685.200 235.800 735.200 236.200 ;
        RECT 685.000 235.600 735.200 235.800 ;
        RECT 764.800 235.800 814.800 236.200 ;
        RECT 764.800 235.600 815.000 235.800 ;
        RECT 685.000 235.200 735.000 235.600 ;
        RECT 684.700 235.000 735.000 235.200 ;
        RECT 765.000 235.200 815.000 235.600 ;
        RECT 765.000 235.000 815.300 235.200 ;
        RECT 684.700 234.600 734.700 235.000 ;
        RECT 684.500 234.400 734.700 234.600 ;
        RECT 765.300 234.600 815.300 235.000 ;
        RECT 765.300 234.400 815.500 234.600 ;
        RECT 684.500 234.000 734.500 234.400 ;
        RECT 684.300 233.800 734.500 234.000 ;
        RECT 765.500 234.000 815.500 234.400 ;
        RECT 765.500 233.800 815.700 234.000 ;
        RECT 684.300 233.400 734.300 233.800 ;
        RECT 684.000 233.200 734.300 233.400 ;
        RECT 765.700 233.400 815.700 233.800 ;
        RECT 765.700 233.200 816.000 233.400 ;
        RECT 684.000 232.800 734.000 233.200 ;
        RECT 683.800 232.600 734.000 232.800 ;
        RECT 766.000 232.800 816.000 233.200 ;
        RECT 766.000 232.600 816.200 232.800 ;
        RECT 683.800 232.200 733.800 232.600 ;
        RECT 683.600 232.000 733.800 232.200 ;
        RECT 766.200 232.200 816.200 232.600 ;
        RECT 766.200 232.000 816.400 232.200 ;
        RECT 683.600 231.600 733.600 232.000 ;
        RECT 683.400 231.400 733.600 231.600 ;
        RECT 766.400 231.600 816.400 232.000 ;
        RECT 766.400 231.400 816.600 231.600 ;
        RECT 683.400 231.000 733.400 231.400 ;
        RECT 683.200 230.800 733.400 231.000 ;
        RECT 766.600 231.000 816.600 231.400 ;
        RECT 766.600 230.800 816.800 231.000 ;
        RECT 683.200 230.400 733.200 230.800 ;
        RECT 682.900 230.200 733.200 230.400 ;
        RECT 766.800 230.400 816.800 230.800 ;
        RECT 766.800 230.200 817.100 230.400 ;
        RECT 682.900 229.800 732.900 230.200 ;
        RECT 682.700 229.600 732.900 229.800 ;
        RECT 767.100 229.800 817.100 230.200 ;
        RECT 767.100 229.600 817.300 229.800 ;
        RECT 682.700 229.200 732.700 229.600 ;
        RECT 682.500 229.000 732.700 229.200 ;
        RECT 767.300 229.200 817.300 229.600 ;
        RECT 767.300 229.000 817.500 229.200 ;
        RECT 682.500 228.600 732.500 229.000 ;
        RECT 682.200 228.400 732.500 228.600 ;
        RECT 767.500 228.600 817.500 229.000 ;
        RECT 767.500 228.400 817.800 228.600 ;
        RECT 682.200 228.000 732.200 228.400 ;
        RECT 682.000 227.800 732.200 228.000 ;
        RECT 767.800 228.000 817.800 228.400 ;
        RECT 767.800 227.800 818.000 228.000 ;
        RECT 682.000 227.400 732.000 227.800 ;
        RECT 681.800 227.200 732.000 227.400 ;
        RECT 768.000 227.400 818.000 227.800 ;
        RECT 768.000 227.200 818.200 227.400 ;
        RECT 681.800 226.800 731.800 227.200 ;
        RECT 681.600 226.600 731.800 226.800 ;
        RECT 768.200 226.800 818.200 227.200 ;
        RECT 768.200 226.600 818.400 226.800 ;
        RECT 681.600 226.200 731.600 226.600 ;
        RECT 681.400 226.000 731.600 226.200 ;
        RECT 768.400 226.200 818.400 226.600 ;
        RECT 768.400 226.000 818.600 226.200 ;
        RECT 681.400 225.600 731.400 226.000 ;
        RECT 681.100 225.400 731.400 225.600 ;
        RECT 768.600 225.600 818.600 226.000 ;
        RECT 768.600 225.400 818.900 225.600 ;
        RECT 681.100 225.000 731.100 225.400 ;
        RECT 680.900 224.800 731.100 225.000 ;
        RECT 768.900 225.000 818.900 225.400 ;
        RECT 768.900 224.800 819.100 225.000 ;
        RECT 680.900 224.400 730.900 224.800 ;
        RECT 680.700 224.200 730.900 224.400 ;
        RECT 769.100 224.400 819.100 224.800 ;
        RECT 769.100 224.200 819.300 224.400 ;
        RECT 680.700 223.800 730.700 224.200 ;
        RECT 680.400 223.600 730.700 223.800 ;
        RECT 769.300 223.800 819.300 224.200 ;
        RECT 769.300 223.600 819.600 223.800 ;
        RECT 680.400 223.200 730.400 223.600 ;
        RECT 680.200 223.000 730.400 223.200 ;
        RECT 769.600 223.200 819.600 223.600 ;
        RECT 769.600 223.000 819.800 223.200 ;
        RECT 680.200 222.600 730.200 223.000 ;
        RECT 680.000 222.400 730.200 222.600 ;
        RECT 769.800 222.600 819.800 223.000 ;
        RECT 769.800 222.400 820.000 222.600 ;
        RECT 680.000 222.000 730.000 222.400 ;
        RECT 679.800 221.800 730.000 222.000 ;
        RECT 770.000 222.000 820.000 222.400 ;
        RECT 770.000 221.800 820.200 222.000 ;
        RECT 679.800 221.400 729.800 221.800 ;
        RECT 679.600 221.200 729.800 221.400 ;
        RECT 770.200 221.400 820.200 221.800 ;
        RECT 770.200 221.200 820.400 221.400 ;
        RECT 679.600 220.800 729.600 221.200 ;
        RECT 679.300 220.600 729.600 220.800 ;
        RECT 770.400 220.800 820.400 221.200 ;
        RECT 770.400 220.600 820.700 220.800 ;
        RECT 679.300 220.200 729.300 220.600 ;
        RECT 679.100 220.000 729.300 220.200 ;
        RECT 770.700 220.200 820.700 220.600 ;
        RECT 770.700 220.000 820.900 220.200 ;
        RECT 679.100 219.600 729.100 220.000 ;
        RECT 678.900 219.400 729.100 219.600 ;
        RECT 770.900 219.600 820.900 220.000 ;
        RECT 770.900 219.400 821.100 219.600 ;
        RECT 678.900 219.000 728.900 219.400 ;
        RECT 678.600 218.800 728.900 219.000 ;
        RECT 771.100 219.000 821.100 219.400 ;
        RECT 771.100 218.800 821.400 219.000 ;
        RECT 678.600 218.400 728.600 218.800 ;
        RECT 678.400 218.200 728.600 218.400 ;
        RECT 771.400 218.400 821.400 218.800 ;
        RECT 771.400 218.200 821.600 218.400 ;
        RECT 678.400 217.800 728.400 218.200 ;
        RECT 678.200 217.600 728.400 217.800 ;
        RECT 771.600 217.800 821.600 218.200 ;
        RECT 771.600 217.600 821.800 217.800 ;
        RECT 678.200 217.200 728.200 217.600 ;
        RECT 678.000 217.000 728.200 217.200 ;
        RECT 771.800 217.200 821.800 217.600 ;
        RECT 771.800 217.000 822.000 217.200 ;
        RECT 678.000 216.600 728.000 217.000 ;
        RECT 677.800 216.400 728.000 216.600 ;
        RECT 772.000 216.600 822.000 217.000 ;
        RECT 772.000 216.400 822.200 216.600 ;
        RECT 677.800 216.000 727.800 216.400 ;
        RECT 677.500 215.800 727.800 216.000 ;
        RECT 772.200 216.000 822.200 216.400 ;
        RECT 772.200 215.800 822.500 216.000 ;
        RECT 677.500 215.400 727.500 215.800 ;
        RECT 677.300 215.200 727.500 215.400 ;
        RECT 772.500 215.400 822.500 215.800 ;
        RECT 772.500 215.200 822.700 215.400 ;
        RECT 677.300 214.800 727.300 215.200 ;
        RECT 677.100 214.600 727.300 214.800 ;
        RECT 772.700 214.800 822.700 215.200 ;
        RECT 772.700 214.600 822.900 214.800 ;
        RECT 677.100 214.200 727.100 214.600 ;
        RECT 676.800 214.000 727.100 214.200 ;
        RECT 772.900 214.200 822.900 214.600 ;
        RECT 772.900 214.000 823.200 214.200 ;
        RECT 676.800 213.600 726.800 214.000 ;
        RECT 676.600 213.400 726.800 213.600 ;
        RECT 773.200 213.600 823.200 214.000 ;
        RECT 773.200 213.400 823.400 213.600 ;
        RECT 676.600 213.000 726.600 213.400 ;
        RECT 676.400 212.800 726.600 213.000 ;
        RECT 773.400 213.000 823.400 213.400 ;
        RECT 773.400 212.800 823.600 213.000 ;
        RECT 676.400 212.400 726.400 212.800 ;
        RECT 676.200 212.200 726.400 212.400 ;
        RECT 773.600 212.400 823.600 212.800 ;
        RECT 773.600 212.200 823.800 212.400 ;
        RECT 676.200 211.800 726.200 212.200 ;
        RECT 676.000 211.600 726.200 211.800 ;
        RECT 773.800 211.800 823.800 212.200 ;
        RECT 773.800 211.600 824.000 211.800 ;
        RECT 676.000 211.200 726.000 211.600 ;
        RECT 675.700 211.000 726.000 211.200 ;
        RECT 774.000 211.200 824.000 211.600 ;
        RECT 774.000 211.000 824.300 211.200 ;
        RECT 675.700 210.600 725.700 211.000 ;
        RECT 675.500 210.400 725.700 210.600 ;
        RECT 774.300 210.600 824.300 211.000 ;
        RECT 774.300 210.400 824.500 210.600 ;
        RECT 675.500 210.000 725.500 210.400 ;
        RECT 675.300 209.800 725.500 210.000 ;
        RECT 774.500 210.000 824.500 210.400 ;
        RECT 774.500 209.800 824.700 210.000 ;
        RECT 675.300 209.400 725.300 209.800 ;
        RECT 675.000 209.200 725.300 209.400 ;
        RECT 774.700 209.400 824.700 209.800 ;
        RECT 774.700 209.200 825.000 209.400 ;
        RECT 675.000 208.800 725.000 209.200 ;
        RECT 674.800 208.600 725.000 208.800 ;
        RECT 775.000 208.800 825.000 209.200 ;
        RECT 775.000 208.600 825.200 208.800 ;
        RECT 674.800 208.200 724.800 208.600 ;
        RECT 674.600 208.000 724.800 208.200 ;
        RECT 775.200 208.200 825.200 208.600 ;
        RECT 775.200 208.000 825.400 208.200 ;
        RECT 674.600 207.600 724.600 208.000 ;
        RECT 674.400 207.400 724.600 207.600 ;
        RECT 775.400 207.600 825.400 208.000 ;
        RECT 775.400 207.400 825.600 207.600 ;
        RECT 674.400 207.000 724.400 207.400 ;
        RECT 674.200 206.800 724.400 207.000 ;
        RECT 775.600 207.000 825.600 207.400 ;
        RECT 775.600 206.800 825.800 207.000 ;
        RECT 674.200 206.400 724.200 206.800 ;
        RECT 673.900 206.200 724.200 206.400 ;
        RECT 775.800 206.400 825.800 206.800 ;
        RECT 775.800 206.200 826.100 206.400 ;
        RECT 673.900 205.800 723.900 206.200 ;
        RECT 673.700 205.600 723.900 205.800 ;
        RECT 776.100 205.800 826.100 206.200 ;
        RECT 776.100 205.600 826.300 205.800 ;
        RECT 673.700 205.200 723.700 205.600 ;
        RECT 673.500 205.000 723.700 205.200 ;
        RECT 776.300 205.200 826.300 205.600 ;
        RECT 776.300 205.000 826.500 205.200 ;
        RECT 673.500 204.600 723.500 205.000 ;
        RECT 673.200 204.400 723.500 204.600 ;
        RECT 776.500 204.600 826.500 205.000 ;
        RECT 776.500 204.400 826.800 204.600 ;
        RECT 673.200 204.000 723.200 204.400 ;
        RECT 673.000 203.800 723.200 204.000 ;
        RECT 776.800 204.000 826.800 204.400 ;
        RECT 776.800 203.800 827.000 204.000 ;
        RECT 673.000 203.400 723.000 203.800 ;
        RECT 672.800 203.200 723.000 203.400 ;
        RECT 777.000 203.400 827.000 203.800 ;
        RECT 777.000 203.200 827.200 203.400 ;
        RECT 672.800 202.800 722.800 203.200 ;
        RECT 672.600 202.600 722.800 202.800 ;
        RECT 777.200 202.800 827.200 203.200 ;
        RECT 777.200 202.600 827.400 202.800 ;
        RECT 672.600 202.200 722.600 202.600 ;
        RECT 672.400 202.000 722.600 202.200 ;
        RECT 777.400 202.200 827.400 202.600 ;
        RECT 777.400 202.000 827.600 202.200 ;
        RECT 672.400 201.600 722.400 202.000 ;
        RECT 672.100 201.400 722.400 201.600 ;
        RECT 777.600 201.600 827.600 202.000 ;
        RECT 777.600 201.400 827.900 201.600 ;
        RECT 672.100 201.000 722.100 201.400 ;
        RECT 671.900 200.800 722.100 201.000 ;
        RECT 777.900 201.000 827.900 201.400 ;
        RECT 777.900 200.800 828.100 201.000 ;
        RECT 671.900 200.400 721.900 200.800 ;
        RECT 671.700 200.200 721.900 200.400 ;
        RECT 778.100 200.400 828.100 200.800 ;
        RECT 778.100 200.200 828.300 200.400 ;
        RECT 671.700 199.800 721.700 200.200 ;
        RECT 671.400 199.600 721.700 199.800 ;
        RECT 778.300 199.800 828.300 200.200 ;
        RECT 778.300 199.600 828.600 199.800 ;
        RECT 671.400 199.200 721.400 199.600 ;
        RECT 671.200 199.000 721.400 199.200 ;
        RECT 778.600 199.200 828.600 199.600 ;
        RECT 778.600 199.000 828.800 199.200 ;
        RECT 671.200 198.600 721.200 199.000 ;
        RECT 671.000 198.400 721.200 198.600 ;
        RECT 778.800 198.600 828.800 199.000 ;
        RECT 778.800 198.400 829.000 198.600 ;
        RECT 671.000 198.000 721.000 198.400 ;
        RECT 670.800 197.800 721.000 198.000 ;
        RECT 779.000 198.000 829.000 198.400 ;
        RECT 779.000 197.800 829.200 198.000 ;
        RECT 670.800 197.400 720.800 197.800 ;
        RECT 670.600 197.200 720.800 197.400 ;
        RECT 779.200 197.400 829.200 197.800 ;
        RECT 779.200 197.200 829.400 197.400 ;
        RECT 670.600 196.800 720.600 197.200 ;
        RECT 670.300 196.600 720.600 196.800 ;
        RECT 779.400 196.800 829.400 197.200 ;
        RECT 779.400 196.600 829.700 196.800 ;
        RECT 670.300 196.200 720.300 196.600 ;
        RECT 670.100 196.000 720.300 196.200 ;
        RECT 779.700 196.200 829.700 196.600 ;
        RECT 779.700 196.000 829.900 196.200 ;
        RECT 670.100 195.600 720.100 196.000 ;
        RECT 669.900 195.400 720.100 195.600 ;
        RECT 779.900 195.600 829.900 196.000 ;
        RECT 779.900 195.400 830.100 195.600 ;
        RECT 669.900 195.000 719.900 195.400 ;
        RECT 669.600 194.800 719.900 195.000 ;
        RECT 780.100 195.000 830.100 195.400 ;
        RECT 780.100 194.800 830.400 195.000 ;
        RECT 669.600 194.400 719.600 194.800 ;
        RECT 669.400 194.200 719.600 194.400 ;
        RECT 780.400 194.400 830.400 194.800 ;
        RECT 780.400 194.200 830.600 194.400 ;
        RECT 669.400 193.800 719.400 194.200 ;
        RECT 669.200 193.600 719.400 193.800 ;
        RECT 780.600 193.800 830.600 194.200 ;
        RECT 780.600 193.600 830.800 193.800 ;
        RECT 669.200 193.200 719.200 193.600 ;
        RECT 669.000 193.000 719.200 193.200 ;
        RECT 780.800 193.200 830.800 193.600 ;
        RECT 780.800 193.000 831.000 193.200 ;
        RECT 669.000 192.600 719.000 193.000 ;
        RECT 668.800 192.400 719.000 192.600 ;
        RECT 781.000 192.600 831.000 193.000 ;
        RECT 781.000 192.400 831.200 192.600 ;
        RECT 668.800 192.000 718.800 192.400 ;
        RECT 668.500 191.800 718.800 192.000 ;
        RECT 781.200 192.000 831.200 192.400 ;
        RECT 781.200 191.800 831.500 192.000 ;
        RECT 668.500 191.400 718.500 191.800 ;
        RECT 668.300 191.200 718.500 191.400 ;
        RECT 781.500 191.400 831.500 191.800 ;
        RECT 781.500 191.200 831.700 191.400 ;
        RECT 668.300 190.800 718.300 191.200 ;
        RECT 668.100 190.600 718.300 190.800 ;
        RECT 781.700 190.800 831.700 191.200 ;
        RECT 781.700 190.600 831.900 190.800 ;
        RECT 668.100 190.200 718.100 190.600 ;
        RECT 667.800 190.000 718.100 190.200 ;
        RECT 781.900 190.200 831.900 190.600 ;
        RECT 781.900 190.000 832.200 190.200 ;
        RECT 667.800 189.600 717.800 190.000 ;
        RECT 667.600 189.400 717.800 189.600 ;
        RECT 782.200 189.600 832.200 190.000 ;
        RECT 782.200 189.400 832.400 189.600 ;
        RECT 667.600 189.000 717.600 189.400 ;
        RECT 667.400 188.800 717.600 189.000 ;
        RECT 782.400 189.000 832.400 189.400 ;
        RECT 782.400 188.800 832.600 189.000 ;
        RECT 667.400 188.400 717.400 188.800 ;
        RECT 667.200 188.200 717.400 188.400 ;
        RECT 782.600 188.400 832.600 188.800 ;
        RECT 782.600 188.200 832.800 188.400 ;
        RECT 667.200 187.800 717.200 188.200 ;
        RECT 667.000 187.600 717.200 187.800 ;
        RECT 782.800 187.800 832.800 188.200 ;
        RECT 782.800 187.600 833.000 187.800 ;
        RECT 667.000 187.200 717.000 187.600 ;
        RECT 666.700 187.000 717.000 187.200 ;
        RECT 783.000 187.200 833.000 187.600 ;
        RECT 783.000 187.000 833.300 187.200 ;
        RECT 666.700 186.600 716.700 187.000 ;
        RECT 666.500 186.400 716.700 186.600 ;
        RECT 783.300 186.600 833.300 187.000 ;
        RECT 783.300 186.400 833.500 186.600 ;
        RECT 666.500 186.000 716.500 186.400 ;
        RECT 666.300 185.800 716.500 186.000 ;
        RECT 783.500 186.000 833.500 186.400 ;
        RECT 783.500 185.800 833.700 186.000 ;
        RECT 666.300 185.400 716.300 185.800 ;
        RECT 666.000 185.200 716.300 185.400 ;
        RECT 783.700 185.400 833.700 185.800 ;
        RECT 783.700 185.200 834.000 185.400 ;
        RECT 666.000 184.800 716.000 185.200 ;
        RECT 665.800 184.600 716.000 184.800 ;
        RECT 784.000 184.800 834.000 185.200 ;
        RECT 784.000 184.600 834.200 184.800 ;
        RECT 665.800 184.200 715.800 184.600 ;
        RECT 665.600 184.000 715.800 184.200 ;
        RECT 784.200 184.200 834.200 184.600 ;
        RECT 784.200 184.000 834.400 184.200 ;
        RECT 665.600 183.600 715.600 184.000 ;
        RECT 665.400 183.400 715.600 183.600 ;
        RECT 784.400 183.600 834.400 184.000 ;
        RECT 784.400 183.400 834.600 183.600 ;
        RECT 665.400 183.000 715.400 183.400 ;
        RECT 665.200 182.800 715.400 183.000 ;
        RECT 784.600 183.000 834.600 183.400 ;
        RECT 784.600 182.800 834.800 183.000 ;
        RECT 665.200 182.400 715.200 182.800 ;
        RECT 664.900 182.200 715.200 182.400 ;
        RECT 784.800 182.400 834.800 182.800 ;
        RECT 784.800 182.200 835.100 182.400 ;
        RECT 664.900 181.800 714.900 182.200 ;
        RECT 664.700 181.600 714.900 181.800 ;
        RECT 785.100 181.800 835.100 182.200 ;
        RECT 785.100 181.600 835.300 181.800 ;
        RECT 664.700 181.200 714.700 181.600 ;
        RECT 664.500 181.000 714.700 181.200 ;
        RECT 785.300 181.200 835.300 181.600 ;
        RECT 785.300 181.000 835.500 181.200 ;
        RECT 664.500 180.600 714.500 181.000 ;
        RECT 664.200 180.400 714.500 180.600 ;
        RECT 785.500 180.600 835.500 181.000 ;
        RECT 785.500 180.400 835.800 180.600 ;
        RECT 664.200 180.000 714.200 180.400 ;
        RECT 664.000 179.800 714.200 180.000 ;
        RECT 785.800 180.000 835.800 180.400 ;
        RECT 785.800 179.800 836.000 180.000 ;
        RECT 664.000 179.400 714.000 179.800 ;
        RECT 663.800 179.200 714.000 179.400 ;
        RECT 786.000 179.400 836.000 179.800 ;
        RECT 786.000 179.200 836.200 179.400 ;
        RECT 663.800 178.800 713.800 179.200 ;
        RECT 663.600 178.600 713.800 178.800 ;
        RECT 786.200 178.800 836.200 179.200 ;
        RECT 786.200 178.600 836.400 178.800 ;
        RECT 663.600 178.200 713.600 178.600 ;
        RECT 663.400 178.000 713.600 178.200 ;
        RECT 786.400 178.200 836.400 178.600 ;
        RECT 786.400 178.000 836.600 178.200 ;
        RECT 663.400 177.600 713.400 178.000 ;
        RECT 663.100 177.400 713.400 177.600 ;
        RECT 786.600 177.600 836.600 178.000 ;
        RECT 786.600 177.400 836.900 177.600 ;
        RECT 663.100 177.000 713.100 177.400 ;
        RECT 662.900 176.800 713.100 177.000 ;
        RECT 786.900 177.000 836.900 177.400 ;
        RECT 786.900 176.800 837.100 177.000 ;
        RECT 662.900 176.400 712.900 176.800 ;
        RECT 662.700 176.200 712.900 176.400 ;
        RECT 787.100 176.400 837.100 176.800 ;
        RECT 787.100 176.200 837.300 176.400 ;
        RECT 662.700 175.800 712.700 176.200 ;
        RECT 662.400 175.600 712.700 175.800 ;
        RECT 787.300 175.800 837.300 176.200 ;
        RECT 787.300 175.600 837.600 175.800 ;
        RECT 662.400 175.200 712.400 175.600 ;
        RECT 662.200 175.000 712.400 175.200 ;
        RECT 787.600 175.200 837.600 175.600 ;
        RECT 787.600 175.000 837.800 175.200 ;
        RECT 662.200 174.600 712.200 175.000 ;
        RECT 662.000 174.400 712.200 174.600 ;
        RECT 787.800 174.600 837.800 175.000 ;
        RECT 787.800 174.400 838.000 174.600 ;
        RECT 662.000 174.000 712.000 174.400 ;
        RECT 661.800 173.800 712.000 174.000 ;
        RECT 788.000 174.000 838.000 174.400 ;
        RECT 788.000 173.800 838.200 174.000 ;
        RECT 661.800 173.400 711.800 173.800 ;
        RECT 661.600 173.200 711.800 173.400 ;
        RECT 788.200 173.400 838.200 173.800 ;
        RECT 788.200 173.200 838.400 173.400 ;
        RECT 661.600 172.800 711.600 173.200 ;
        RECT 661.300 172.600 711.600 172.800 ;
        RECT 788.400 172.800 838.400 173.200 ;
        RECT 788.400 172.600 838.700 172.800 ;
        RECT 661.300 172.200 711.300 172.600 ;
        RECT 661.100 172.000 711.300 172.200 ;
        RECT 788.700 172.200 838.700 172.600 ;
        RECT 788.700 172.000 838.900 172.200 ;
        RECT 661.100 171.600 711.100 172.000 ;
        RECT 660.900 171.400 711.100 171.600 ;
        RECT 788.900 171.600 838.900 172.000 ;
        RECT 788.900 171.400 839.100 171.600 ;
        RECT 660.900 171.000 710.900 171.400 ;
        RECT 660.600 170.800 710.900 171.000 ;
        RECT 789.100 171.000 839.100 171.400 ;
        RECT 789.100 170.800 839.400 171.000 ;
        RECT 660.600 170.400 710.600 170.800 ;
        RECT 660.400 170.200 710.600 170.400 ;
        RECT 789.400 170.400 839.400 170.800 ;
        RECT 789.400 170.200 839.600 170.400 ;
        RECT 660.400 169.800 710.400 170.200 ;
        RECT 660.200 169.600 710.400 169.800 ;
        RECT 789.600 169.800 839.600 170.200 ;
        RECT 789.600 169.600 839.800 169.800 ;
        RECT 660.200 169.200 710.200 169.600 ;
        RECT 660.000 169.000 710.200 169.200 ;
        RECT 789.800 169.200 839.800 169.600 ;
        RECT 789.800 169.000 840.000 169.200 ;
        RECT 660.000 168.600 710.000 169.000 ;
        RECT 659.800 168.400 710.000 168.600 ;
        RECT 790.000 168.600 840.000 169.000 ;
        RECT 790.000 168.400 840.200 168.600 ;
        RECT 659.800 168.000 709.800 168.400 ;
        RECT 659.500 167.800 709.800 168.000 ;
        RECT 790.200 168.000 840.200 168.400 ;
        RECT 790.200 167.800 840.500 168.000 ;
        RECT 659.500 167.400 709.500 167.800 ;
        RECT 659.300 167.200 709.500 167.400 ;
        RECT 790.500 167.400 840.500 167.800 ;
        RECT 790.500 167.200 840.700 167.400 ;
        RECT 659.300 166.800 709.300 167.200 ;
        RECT 659.100 166.600 709.300 166.800 ;
        RECT 790.700 166.800 840.700 167.200 ;
        RECT 790.700 166.600 840.900 166.800 ;
        RECT 659.100 166.200 709.100 166.600 ;
        RECT 658.800 166.000 709.100 166.200 ;
        RECT 790.900 166.200 840.900 166.600 ;
        RECT 790.900 166.000 841.200 166.200 ;
        RECT 658.800 165.600 708.800 166.000 ;
        RECT 658.600 165.400 708.800 165.600 ;
        RECT 791.200 165.600 841.200 166.000 ;
        RECT 791.200 165.400 841.400 165.600 ;
        RECT 658.600 165.000 708.600 165.400 ;
        RECT 658.400 164.800 708.600 165.000 ;
        RECT 791.400 165.000 841.400 165.400 ;
        RECT 791.400 164.800 841.600 165.000 ;
        RECT 658.400 164.400 708.400 164.800 ;
        RECT 658.200 164.200 708.400 164.400 ;
        RECT 791.600 164.400 841.600 164.800 ;
        RECT 791.600 164.200 841.800 164.400 ;
        RECT 658.200 163.800 708.200 164.200 ;
        RECT 658.000 163.600 708.200 163.800 ;
        RECT 791.800 163.800 841.800 164.200 ;
        RECT 791.800 163.600 842.000 163.800 ;
        RECT 658.000 163.200 708.000 163.600 ;
        RECT 657.700 163.000 708.000 163.200 ;
        RECT 792.000 163.200 842.000 163.600 ;
        RECT 792.000 163.000 842.300 163.200 ;
        RECT 657.700 162.600 707.700 163.000 ;
        RECT 657.500 162.400 707.700 162.600 ;
        RECT 792.300 162.600 842.300 163.000 ;
        RECT 792.300 162.400 842.500 162.600 ;
        RECT 657.500 162.000 707.500 162.400 ;
        RECT 792.500 162.000 842.500 162.400 ;
        RECT 657.300 161.400 842.700 162.000 ;
        RECT 657.000 160.800 843.000 161.400 ;
        RECT 656.800 160.200 843.200 160.800 ;
        RECT 656.600 159.600 843.400 160.200 ;
        RECT 656.400 159.000 843.600 159.600 ;
        RECT 656.200 158.400 843.800 159.000 ;
        RECT 655.900 157.800 844.100 158.400 ;
        RECT 655.700 157.200 844.300 157.800 ;
        RECT 655.500 156.600 844.500 157.200 ;
        RECT 655.200 156.000 844.800 156.600 ;
        RECT 655.000 155.400 845.000 156.000 ;
        RECT 654.800 154.800 845.200 155.400 ;
        RECT 654.600 154.200 845.400 154.800 ;
        RECT 654.400 153.600 845.600 154.200 ;
        RECT 654.100 153.000 845.900 153.600 ;
        RECT 653.900 152.400 846.100 153.000 ;
        RECT 653.700 151.800 846.300 152.400 ;
        RECT 653.400 151.200 846.600 151.800 ;
        RECT 653.200 150.600 846.800 151.200 ;
        RECT 653.000 150.000 847.000 150.600 ;
        RECT 652.800 149.400 847.200 150.000 ;
        RECT 652.600 148.800 847.400 149.400 ;
        RECT 652.300 148.200 847.700 148.800 ;
        RECT 652.100 147.600 847.900 148.200 ;
        RECT 651.900 147.000 848.100 147.600 ;
        RECT 651.600 146.400 848.400 147.000 ;
        RECT 651.400 145.800 848.600 146.400 ;
        RECT 651.200 145.200 848.800 145.800 ;
        RECT 651.000 144.600 849.000 145.200 ;
        RECT 650.800 144.000 849.200 144.600 ;
        RECT 650.500 143.400 849.500 144.000 ;
        RECT 650.300 142.800 849.700 143.400 ;
        RECT 650.100 142.200 849.900 142.800 ;
        RECT 649.800 141.600 850.200 142.200 ;
        RECT 649.600 141.000 850.400 141.600 ;
        RECT 649.400 140.400 850.600 141.000 ;
        RECT 649.200 139.800 850.800 140.400 ;
        RECT 649.000 139.200 851.000 139.800 ;
        RECT 648.700 138.600 851.300 139.200 ;
        RECT 648.500 138.000 851.500 138.600 ;
        RECT 648.300 137.400 851.700 138.000 ;
        RECT 648.000 136.800 852.000 137.400 ;
        RECT 647.800 136.200 852.200 136.800 ;
        RECT 647.600 135.600 852.400 136.200 ;
        RECT 647.400 135.000 852.600 135.600 ;
        RECT 647.200 134.400 852.800 135.000 ;
        RECT 646.900 133.800 853.100 134.400 ;
        RECT 646.700 133.200 853.300 133.800 ;
        RECT 646.500 132.600 853.500 133.200 ;
        RECT 646.200 132.000 853.800 132.600 ;
        RECT 646.000 131.400 854.000 132.000 ;
        RECT 645.800 130.800 854.200 131.400 ;
        RECT 645.600 130.200 854.400 130.800 ;
        RECT 645.400 129.600 854.600 130.200 ;
        RECT 645.100 129.000 854.900 129.600 ;
        RECT 644.900 128.400 855.100 129.000 ;
        RECT 644.700 127.800 855.300 128.400 ;
        RECT 644.400 127.200 855.600 127.800 ;
        RECT 644.200 126.600 855.800 127.200 ;
        RECT 644.000 126.000 856.000 126.600 ;
        RECT 643.800 125.400 856.200 126.000 ;
        RECT 643.600 124.800 856.400 125.400 ;
        RECT 643.300 124.200 856.700 124.800 ;
        RECT 643.100 123.600 856.900 124.200 ;
        RECT 642.900 123.000 857.100 123.600 ;
        RECT 642.600 122.400 857.400 123.000 ;
        RECT 642.400 122.200 857.600 122.400 ;
        RECT 642.400 121.800 692.400 122.200 ;
        RECT 642.200 121.600 692.400 121.800 ;
        RECT 807.600 121.800 857.600 122.200 ;
        RECT 807.600 121.600 857.800 121.800 ;
        RECT 642.200 121.200 692.200 121.600 ;
        RECT 642.000 121.000 692.200 121.200 ;
        RECT 807.800 121.200 857.800 121.600 ;
        RECT 807.800 121.000 858.000 121.200 ;
        RECT 642.000 120.600 692.000 121.000 ;
        RECT 641.800 120.400 692.000 120.600 ;
        RECT 808.000 120.600 858.000 121.000 ;
        RECT 808.000 120.400 858.200 120.600 ;
        RECT 641.800 120.000 691.800 120.400 ;
        RECT 641.500 119.800 691.800 120.000 ;
        RECT 808.200 120.000 858.200 120.400 ;
        RECT 808.200 119.800 858.500 120.000 ;
        RECT 641.500 119.400 691.500 119.800 ;
        RECT 641.300 119.200 691.500 119.400 ;
        RECT 808.500 119.400 858.500 119.800 ;
        RECT 808.500 119.200 858.700 119.400 ;
        RECT 641.300 118.800 691.300 119.200 ;
        RECT 641.100 118.600 691.300 118.800 ;
        RECT 808.700 118.800 858.700 119.200 ;
        RECT 808.700 118.600 858.900 118.800 ;
        RECT 641.100 118.200 691.100 118.600 ;
        RECT 640.800 118.000 691.100 118.200 ;
        RECT 808.900 118.200 858.900 118.600 ;
        RECT 808.900 118.000 859.200 118.200 ;
        RECT 640.800 117.600 690.800 118.000 ;
        RECT 640.600 117.400 690.800 117.600 ;
        RECT 809.200 117.600 859.200 118.000 ;
        RECT 809.200 117.400 859.400 117.600 ;
        RECT 640.600 117.000 690.600 117.400 ;
        RECT 640.400 116.800 690.600 117.000 ;
        RECT 809.400 117.000 859.400 117.400 ;
        RECT 809.400 116.800 859.600 117.000 ;
        RECT 640.400 116.400 690.400 116.800 ;
        RECT 640.200 116.200 690.400 116.400 ;
        RECT 809.600 116.400 859.600 116.800 ;
        RECT 809.600 116.200 859.800 116.400 ;
        RECT 640.200 115.800 690.200 116.200 ;
        RECT 640.000 115.600 690.200 115.800 ;
        RECT 809.800 115.800 859.800 116.200 ;
        RECT 809.800 115.600 860.000 115.800 ;
        RECT 640.000 115.200 690.000 115.600 ;
        RECT 639.700 115.000 690.000 115.200 ;
        RECT 810.000 115.200 860.000 115.600 ;
        RECT 810.000 115.000 860.300 115.200 ;
        RECT 639.700 114.600 689.700 115.000 ;
        RECT 639.500 114.400 689.700 114.600 ;
        RECT 810.300 114.600 860.300 115.000 ;
        RECT 810.300 114.400 860.500 114.600 ;
        RECT 639.500 114.000 689.500 114.400 ;
        RECT 639.300 113.800 689.500 114.000 ;
        RECT 810.500 114.000 860.500 114.400 ;
        RECT 810.500 113.800 860.700 114.000 ;
        RECT 639.300 113.400 689.300 113.800 ;
        RECT 639.000 113.200 689.300 113.400 ;
        RECT 810.700 113.400 860.700 113.800 ;
        RECT 810.700 113.200 861.000 113.400 ;
        RECT 639.000 112.800 689.000 113.200 ;
        RECT 638.800 112.600 689.000 112.800 ;
        RECT 811.000 112.800 861.000 113.200 ;
        RECT 811.000 112.600 861.200 112.800 ;
        RECT 638.800 112.200 688.800 112.600 ;
        RECT 638.600 112.000 688.800 112.200 ;
        RECT 811.200 112.200 861.200 112.600 ;
        RECT 811.200 112.000 861.400 112.200 ;
        RECT 638.600 111.600 688.600 112.000 ;
        RECT 638.400 111.400 688.600 111.600 ;
        RECT 811.400 111.600 861.400 112.000 ;
        RECT 811.400 111.400 861.600 111.600 ;
        RECT 638.400 111.000 688.400 111.400 ;
        RECT 638.200 110.800 688.400 111.000 ;
        RECT 811.600 111.000 861.600 111.400 ;
        RECT 811.600 110.800 861.800 111.000 ;
        RECT 638.200 110.400 688.200 110.800 ;
        RECT 637.900 110.200 688.200 110.400 ;
        RECT 811.800 110.400 861.800 110.800 ;
        RECT 811.800 110.200 862.100 110.400 ;
        RECT 637.900 109.800 687.900 110.200 ;
        RECT 637.700 109.600 687.900 109.800 ;
        RECT 812.100 109.800 862.100 110.200 ;
        RECT 812.100 109.600 862.300 109.800 ;
        RECT 637.700 109.200 687.700 109.600 ;
        RECT 637.500 109.000 687.700 109.200 ;
        RECT 812.300 109.200 862.300 109.600 ;
        RECT 812.300 109.000 862.500 109.200 ;
        RECT 637.500 108.600 687.500 109.000 ;
        RECT 637.200 108.400 687.500 108.600 ;
        RECT 812.500 108.600 862.500 109.000 ;
        RECT 812.500 108.400 862.800 108.600 ;
        RECT 637.200 108.000 687.200 108.400 ;
        RECT 637.000 107.800 687.200 108.000 ;
        RECT 812.800 108.000 862.800 108.400 ;
        RECT 812.800 107.800 863.000 108.000 ;
        RECT 637.000 107.400 687.000 107.800 ;
        RECT 636.800 107.200 687.000 107.400 ;
        RECT 813.000 107.400 863.000 107.800 ;
        RECT 813.000 107.200 863.200 107.400 ;
        RECT 636.800 106.800 686.800 107.200 ;
        RECT 636.600 106.600 686.800 106.800 ;
        RECT 813.200 106.800 863.200 107.200 ;
        RECT 813.200 106.600 863.400 106.800 ;
        RECT 636.600 106.200 686.600 106.600 ;
        RECT 636.400 106.000 686.600 106.200 ;
        RECT 813.400 106.200 863.400 106.600 ;
        RECT 813.400 106.000 863.600 106.200 ;
        RECT 636.400 105.600 686.400 106.000 ;
        RECT 636.100 105.400 686.400 105.600 ;
        RECT 813.600 105.600 863.600 106.000 ;
        RECT 813.600 105.400 863.900 105.600 ;
        RECT 636.100 105.000 686.100 105.400 ;
        RECT 635.900 104.800 686.100 105.000 ;
        RECT 813.900 105.000 863.900 105.400 ;
        RECT 813.900 104.800 864.100 105.000 ;
        RECT 635.900 104.400 685.900 104.800 ;
        RECT 635.700 104.200 685.900 104.400 ;
        RECT 814.100 104.400 864.100 104.800 ;
        RECT 814.100 104.200 864.300 104.400 ;
        RECT 635.700 103.800 685.700 104.200 ;
        RECT 635.400 103.600 685.700 103.800 ;
        RECT 814.300 103.800 864.300 104.200 ;
        RECT 814.300 103.600 864.600 103.800 ;
        RECT 635.400 103.200 685.400 103.600 ;
        RECT 635.200 103.000 685.400 103.200 ;
        RECT 814.600 103.200 864.600 103.600 ;
        RECT 814.600 103.000 864.800 103.200 ;
        RECT 635.200 102.600 685.200 103.000 ;
        RECT 635.000 102.400 685.200 102.600 ;
        RECT 814.800 102.600 864.800 103.000 ;
        RECT 814.800 102.400 865.000 102.600 ;
        RECT 635.000 102.000 685.000 102.400 ;
        RECT 634.800 101.800 685.000 102.000 ;
        RECT 815.000 102.000 865.000 102.400 ;
        RECT 815.000 101.800 865.200 102.000 ;
        RECT 634.800 101.400 684.800 101.800 ;
        RECT 634.600 101.200 684.800 101.400 ;
        RECT 815.200 101.400 865.200 101.800 ;
        RECT 815.200 101.200 865.400 101.400 ;
        RECT 634.600 100.800 684.600 101.200 ;
        RECT 634.300 100.600 684.600 100.800 ;
        RECT 815.400 100.800 865.400 101.200 ;
        RECT 815.400 100.600 865.700 100.800 ;
        RECT 634.300 100.200 684.300 100.600 ;
        RECT 634.100 100.000 684.300 100.200 ;
        RECT 815.700 100.200 865.700 100.600 ;
        RECT 815.700 100.000 865.900 100.200 ;
        RECT 634.100 99.600 684.100 100.000 ;
        RECT 633.900 99.400 684.100 99.600 ;
        RECT 815.900 99.600 865.900 100.000 ;
        RECT 815.900 99.400 866.100 99.600 ;
        RECT 633.900 99.000 683.900 99.400 ;
        RECT 633.600 98.800 683.900 99.000 ;
        RECT 816.100 99.000 866.100 99.400 ;
        RECT 816.100 98.800 866.400 99.000 ;
        RECT 633.600 98.400 683.600 98.800 ;
        RECT 633.400 98.200 683.600 98.400 ;
        RECT 816.400 98.400 866.400 98.800 ;
        RECT 816.400 98.200 866.600 98.400 ;
        RECT 633.400 97.800 683.400 98.200 ;
        RECT 633.200 97.600 683.400 97.800 ;
        RECT 816.600 97.800 866.600 98.200 ;
        RECT 816.600 97.600 866.800 97.800 ;
        RECT 633.200 97.200 683.200 97.600 ;
        RECT 633.000 97.000 683.200 97.200 ;
        RECT 816.800 97.200 866.800 97.600 ;
        RECT 816.800 97.000 867.000 97.200 ;
        RECT 633.000 96.600 683.000 97.000 ;
        RECT 632.800 96.400 683.000 96.600 ;
        RECT 817.000 96.600 867.000 97.000 ;
        RECT 817.000 96.400 867.200 96.600 ;
        RECT 632.800 96.000 682.800 96.400 ;
        RECT 632.500 95.800 682.800 96.000 ;
        RECT 817.200 96.000 867.200 96.400 ;
        RECT 817.200 95.800 867.500 96.000 ;
        RECT 632.500 95.400 682.500 95.800 ;
        RECT 632.300 95.200 682.500 95.400 ;
        RECT 817.500 95.400 867.500 95.800 ;
        RECT 817.500 95.200 867.700 95.400 ;
        RECT 632.300 94.800 682.300 95.200 ;
        RECT 632.100 94.600 682.300 94.800 ;
        RECT 817.700 94.800 867.700 95.200 ;
        RECT 817.700 94.600 867.900 94.800 ;
        RECT 632.100 94.200 682.100 94.600 ;
        RECT 631.800 94.000 682.100 94.200 ;
        RECT 817.900 94.200 867.900 94.600 ;
        RECT 817.900 94.000 868.200 94.200 ;
        RECT 631.800 93.600 681.800 94.000 ;
        RECT 631.600 93.400 681.800 93.600 ;
        RECT 818.200 93.600 868.200 94.000 ;
        RECT 818.200 93.400 868.400 93.600 ;
        RECT 631.600 93.000 681.600 93.400 ;
        RECT 631.400 92.800 681.600 93.000 ;
        RECT 818.400 93.000 868.400 93.400 ;
        RECT 818.400 92.800 868.600 93.000 ;
        RECT 631.400 92.400 681.400 92.800 ;
        RECT 631.200 92.200 681.400 92.400 ;
        RECT 818.600 92.400 868.600 92.800 ;
        RECT 818.600 92.200 868.800 92.400 ;
        RECT 631.200 91.800 681.200 92.200 ;
        RECT 631.000 91.600 681.200 91.800 ;
        RECT 818.800 91.800 868.800 92.200 ;
        RECT 818.800 91.600 869.000 91.800 ;
        RECT 631.000 91.200 681.000 91.600 ;
        RECT 630.700 91.000 681.000 91.200 ;
        RECT 819.000 91.200 869.000 91.600 ;
        RECT 819.000 91.000 869.300 91.200 ;
        RECT 630.700 90.600 680.700 91.000 ;
        RECT 630.500 90.400 680.700 90.600 ;
        RECT 819.300 90.600 869.300 91.000 ;
        RECT 819.300 90.400 869.500 90.600 ;
        RECT 630.500 90.000 680.500 90.400 ;
        RECT 630.300 89.800 680.500 90.000 ;
        RECT 819.500 90.000 869.500 90.400 ;
        RECT 819.500 89.800 869.700 90.000 ;
        RECT 630.300 89.400 680.300 89.800 ;
        RECT 630.000 89.200 680.300 89.400 ;
        RECT 819.700 89.400 869.700 89.800 ;
        RECT 819.700 89.200 870.000 89.400 ;
        RECT 630.000 88.800 680.000 89.200 ;
        RECT 629.800 88.600 680.000 88.800 ;
        RECT 820.000 88.800 870.000 89.200 ;
        RECT 820.000 88.600 870.200 88.800 ;
        RECT 629.800 88.200 679.800 88.600 ;
        RECT 629.600 88.000 679.800 88.200 ;
        RECT 820.200 88.200 870.200 88.600 ;
        RECT 820.200 88.000 870.400 88.200 ;
        RECT 629.600 87.600 679.600 88.000 ;
        RECT 629.400 87.400 679.600 87.600 ;
        RECT 820.400 87.600 870.400 88.000 ;
        RECT 820.400 87.400 870.600 87.600 ;
        RECT 629.400 87.000 679.400 87.400 ;
        RECT 629.200 86.800 679.400 87.000 ;
        RECT 820.600 87.000 870.600 87.400 ;
        RECT 820.600 86.800 870.800 87.000 ;
        RECT 629.200 86.400 679.200 86.800 ;
        RECT 628.900 86.200 679.200 86.400 ;
        RECT 820.800 86.400 870.800 86.800 ;
        RECT 820.800 86.200 871.100 86.400 ;
        RECT 628.900 85.800 678.900 86.200 ;
        RECT 628.700 85.600 678.900 85.800 ;
        RECT 821.100 85.800 871.100 86.200 ;
        RECT 821.100 85.600 871.300 85.800 ;
        RECT 628.700 85.200 678.700 85.600 ;
        RECT 628.500 85.000 678.700 85.200 ;
        RECT 821.300 85.200 871.300 85.600 ;
        RECT 821.300 85.000 871.500 85.200 ;
        RECT 628.500 84.600 678.500 85.000 ;
        RECT 628.200 84.400 678.500 84.600 ;
        RECT 821.500 84.600 871.500 85.000 ;
        RECT 821.500 84.400 871.800 84.600 ;
        RECT 628.200 84.000 678.200 84.400 ;
        RECT 628.000 83.800 678.200 84.000 ;
        RECT 821.800 84.000 871.800 84.400 ;
        RECT 821.800 83.800 872.000 84.000 ;
        RECT 628.000 83.400 678.000 83.800 ;
        RECT 627.800 83.200 678.000 83.400 ;
        RECT 822.000 83.400 872.000 83.800 ;
        RECT 822.000 83.200 872.200 83.400 ;
        RECT 627.800 82.800 677.800 83.200 ;
        RECT 627.600 82.600 677.800 82.800 ;
        RECT 822.200 82.800 872.200 83.200 ;
        RECT 822.200 82.600 872.400 82.800 ;
        RECT 627.600 82.200 677.600 82.600 ;
        RECT 627.400 82.000 677.600 82.200 ;
        RECT 822.400 82.200 872.400 82.600 ;
        RECT 822.400 82.000 872.600 82.200 ;
        RECT 627.400 81.600 677.400 82.000 ;
        RECT 627.100 81.400 677.400 81.600 ;
        RECT 822.600 81.600 872.600 82.000 ;
        RECT 822.600 81.400 872.900 81.600 ;
        RECT 627.100 81.000 677.100 81.400 ;
        RECT 626.900 80.800 677.100 81.000 ;
        RECT 822.900 81.000 872.900 81.400 ;
        RECT 822.900 80.800 873.100 81.000 ;
        RECT 626.900 80.400 676.900 80.800 ;
        RECT 626.700 80.200 676.900 80.400 ;
        RECT 823.100 80.400 873.100 80.800 ;
        RECT 823.100 80.200 873.300 80.400 ;
        RECT 626.700 79.800 676.700 80.200 ;
        RECT 626.400 79.600 676.700 79.800 ;
        RECT 823.300 79.800 873.300 80.200 ;
        RECT 823.300 79.600 873.600 79.800 ;
        RECT 626.400 79.200 676.400 79.600 ;
        RECT 626.200 79.000 676.400 79.200 ;
        RECT 823.600 79.200 873.600 79.600 ;
        RECT 823.600 79.000 873.800 79.200 ;
        RECT 626.200 78.600 676.200 79.000 ;
        RECT 626.000 78.400 676.200 78.600 ;
        RECT 823.800 78.600 873.800 79.000 ;
        RECT 823.800 78.400 874.000 78.600 ;
        RECT 626.000 78.000 676.000 78.400 ;
        RECT 625.800 77.800 676.000 78.000 ;
        RECT 824.000 78.000 874.000 78.400 ;
        RECT 824.000 77.800 874.200 78.000 ;
        RECT 625.800 77.400 675.800 77.800 ;
        RECT 625.600 77.200 675.800 77.400 ;
        RECT 824.200 77.400 874.200 77.800 ;
        RECT 824.200 77.200 874.400 77.400 ;
        RECT 625.600 76.800 675.600 77.200 ;
        RECT 625.300 76.600 675.600 76.800 ;
        RECT 824.400 76.800 874.400 77.200 ;
        RECT 824.400 76.600 874.700 76.800 ;
        RECT 625.300 76.200 675.300 76.600 ;
        RECT 625.100 76.000 675.300 76.200 ;
        RECT 824.700 76.200 874.700 76.600 ;
        RECT 824.700 76.000 874.900 76.200 ;
        RECT 625.100 75.600 675.100 76.000 ;
        RECT 624.900 75.400 675.100 75.600 ;
        RECT 824.900 75.600 874.900 76.000 ;
        RECT 824.900 75.400 875.100 75.600 ;
        RECT 624.900 75.000 674.900 75.400 ;
        RECT 624.600 74.800 674.900 75.000 ;
        RECT 825.100 75.000 875.100 75.400 ;
        RECT 825.100 74.800 875.400 75.000 ;
        RECT 624.600 74.400 674.600 74.800 ;
        RECT 624.400 74.200 674.600 74.400 ;
        RECT 825.400 74.400 875.400 74.800 ;
        RECT 825.400 74.200 875.600 74.400 ;
        RECT 624.400 73.800 674.400 74.200 ;
        RECT 624.200 73.600 674.400 73.800 ;
        RECT 825.600 73.800 875.600 74.200 ;
        RECT 825.600 73.600 875.800 73.800 ;
        RECT 624.200 73.200 674.200 73.600 ;
        RECT 624.000 73.000 674.200 73.200 ;
        RECT 825.800 73.200 875.800 73.600 ;
        RECT 825.800 73.000 876.000 73.200 ;
        RECT 624.000 72.600 674.000 73.000 ;
        RECT 623.800 72.400 674.000 72.600 ;
        RECT 826.000 72.600 876.000 73.000 ;
        RECT 826.000 72.400 876.200 72.600 ;
        RECT 623.800 72.000 673.800 72.400 ;
        RECT 623.500 71.800 673.800 72.000 ;
        RECT 826.200 72.000 876.200 72.400 ;
        RECT 826.200 71.800 876.500 72.000 ;
        RECT 623.500 71.400 673.500 71.800 ;
        RECT 623.300 71.200 673.500 71.400 ;
        RECT 826.500 71.400 876.500 71.800 ;
        RECT 826.500 71.200 876.700 71.400 ;
        RECT 623.300 70.800 673.300 71.200 ;
        RECT 623.100 70.600 673.300 70.800 ;
        RECT 826.700 70.800 876.700 71.200 ;
        RECT 826.700 70.600 876.900 70.800 ;
        RECT 623.100 70.200 673.100 70.600 ;
        RECT 622.800 70.000 673.100 70.200 ;
        RECT 826.900 70.200 876.900 70.600 ;
        RECT 826.900 70.000 877.200 70.200 ;
        RECT 622.800 69.600 672.800 70.000 ;
        RECT 622.600 69.400 672.800 69.600 ;
        RECT 827.200 69.600 877.200 70.000 ;
        RECT 827.200 69.400 877.400 69.600 ;
        RECT 622.600 69.000 672.600 69.400 ;
        RECT 622.400 68.800 672.600 69.000 ;
        RECT 827.400 69.000 877.400 69.400 ;
        RECT 827.400 68.800 877.600 69.000 ;
        RECT 622.400 68.400 672.400 68.800 ;
        RECT 622.200 68.200 672.400 68.400 ;
        RECT 827.600 68.400 877.600 68.800 ;
        RECT 827.600 68.200 877.800 68.400 ;
        RECT 622.200 67.800 672.200 68.200 ;
        RECT 622.000 67.600 672.200 67.800 ;
        RECT 827.800 67.800 877.800 68.200 ;
        RECT 827.800 67.600 878.000 67.800 ;
        RECT 622.000 67.200 672.000 67.600 ;
        RECT 621.700 67.000 672.000 67.200 ;
        RECT 828.000 67.200 878.000 67.600 ;
        RECT 828.000 67.000 878.300 67.200 ;
        RECT 621.700 66.600 671.700 67.000 ;
        RECT 621.500 66.400 671.700 66.600 ;
        RECT 828.300 66.600 878.300 67.000 ;
        RECT 828.300 66.400 878.500 66.600 ;
        RECT 621.500 66.000 671.500 66.400 ;
        RECT 621.300 65.800 671.500 66.000 ;
        RECT 828.500 66.000 878.500 66.400 ;
        RECT 828.500 65.800 878.700 66.000 ;
        RECT 621.300 65.400 671.300 65.800 ;
        RECT 621.000 65.200 671.300 65.400 ;
        RECT 828.700 65.400 878.700 65.800 ;
        RECT 828.700 65.200 879.000 65.400 ;
        RECT 621.000 64.800 671.000 65.200 ;
        RECT 620.800 64.600 671.000 64.800 ;
        RECT 829.000 64.800 879.000 65.200 ;
        RECT 829.000 64.600 879.200 64.800 ;
        RECT 620.800 64.200 670.800 64.600 ;
        RECT 620.600 64.000 670.800 64.200 ;
        RECT 829.200 64.200 879.200 64.600 ;
        RECT 829.200 64.000 879.400 64.200 ;
        RECT 620.600 63.600 670.600 64.000 ;
        RECT 620.400 63.400 670.600 63.600 ;
        RECT 829.400 63.600 879.400 64.000 ;
        RECT 829.400 63.400 879.600 63.600 ;
        RECT 620.400 63.000 670.400 63.400 ;
        RECT 620.200 62.800 670.400 63.000 ;
        RECT 829.600 63.000 879.600 63.400 ;
        RECT 829.600 62.800 879.800 63.000 ;
        RECT 620.200 62.400 670.200 62.800 ;
        RECT 619.900 62.200 670.200 62.400 ;
        RECT 829.800 62.400 879.800 62.800 ;
        RECT 829.800 62.200 880.100 62.400 ;
        RECT 619.900 61.800 669.900 62.200 ;
        RECT 619.700 61.600 669.900 61.800 ;
        RECT 830.100 61.800 880.100 62.200 ;
        RECT 830.100 61.600 880.300 61.800 ;
        RECT 619.700 61.200 669.700 61.600 ;
        RECT 619.500 61.000 669.700 61.200 ;
        RECT 830.300 61.200 880.300 61.600 ;
        RECT 830.300 61.000 880.500 61.200 ;
        RECT 619.500 60.600 669.500 61.000 ;
        RECT 619.200 60.400 669.500 60.600 ;
        RECT 830.500 60.600 880.500 61.000 ;
        RECT 830.500 60.400 880.800 60.600 ;
        RECT 619.200 60.000 669.200 60.400 ;
        RECT 619.000 59.800 669.200 60.000 ;
        RECT 830.800 60.000 880.800 60.400 ;
        RECT 830.800 59.800 881.000 60.000 ;
        RECT 619.000 59.400 669.000 59.800 ;
        RECT 618.800 59.200 669.000 59.400 ;
        RECT 831.000 59.400 881.000 59.800 ;
        RECT 831.000 59.200 881.200 59.400 ;
        RECT 618.800 58.800 668.800 59.200 ;
        RECT 618.600 58.600 668.800 58.800 ;
        RECT 831.200 58.800 881.200 59.200 ;
        RECT 831.200 58.600 881.400 58.800 ;
        RECT 618.600 58.200 668.600 58.600 ;
        RECT 618.400 58.000 668.600 58.200 ;
        RECT 831.400 58.200 881.400 58.600 ;
        RECT 831.400 58.000 881.600 58.200 ;
        RECT 618.400 57.600 668.400 58.000 ;
        RECT 618.100 57.400 668.400 57.600 ;
        RECT 831.600 57.600 881.600 58.000 ;
        RECT 831.600 57.400 881.900 57.600 ;
        RECT 618.100 57.000 668.100 57.400 ;
        RECT 617.900 56.800 668.100 57.000 ;
        RECT 831.900 57.000 881.900 57.400 ;
        RECT 831.900 56.800 882.100 57.000 ;
        RECT 617.900 56.400 667.900 56.800 ;
        RECT 617.700 56.200 667.900 56.400 ;
        RECT 832.100 56.400 882.100 56.800 ;
        RECT 832.100 56.200 882.300 56.400 ;
        RECT 617.700 55.800 667.700 56.200 ;
        RECT 617.400 55.600 667.700 55.800 ;
        RECT 832.300 55.800 882.300 56.200 ;
        RECT 832.300 55.600 882.600 55.800 ;
        RECT 617.400 55.200 667.400 55.600 ;
        RECT 617.200 55.000 667.400 55.200 ;
        RECT 832.600 55.200 882.600 55.600 ;
        RECT 832.600 55.000 882.800 55.200 ;
        RECT 617.200 54.600 667.200 55.000 ;
        RECT 617.000 54.400 667.200 54.600 ;
        RECT 832.800 54.600 882.800 55.000 ;
        RECT 832.800 54.400 883.000 54.600 ;
        RECT 617.000 54.000 667.000 54.400 ;
        RECT 616.800 53.800 667.000 54.000 ;
        RECT 833.000 54.000 883.000 54.400 ;
        RECT 833.000 53.800 883.200 54.000 ;
        RECT 616.800 53.400 666.800 53.800 ;
        RECT 616.600 53.200 666.800 53.400 ;
        RECT 833.200 53.400 883.200 53.800 ;
        RECT 833.200 53.200 883.400 53.400 ;
        RECT 616.600 52.800 666.600 53.200 ;
        RECT 616.300 52.600 666.600 52.800 ;
        RECT 833.400 52.800 883.400 53.200 ;
        RECT 833.400 52.600 883.700 52.800 ;
        RECT 616.300 52.200 666.300 52.600 ;
        RECT 616.100 52.000 666.300 52.200 ;
        RECT 833.700 52.200 883.700 52.600 ;
        RECT 833.700 52.000 883.900 52.200 ;
        RECT 616.100 51.600 666.100 52.000 ;
        RECT 615.900 51.400 666.100 51.600 ;
        RECT 833.900 51.600 883.900 52.000 ;
        RECT 833.900 51.400 884.100 51.600 ;
        RECT 615.900 51.000 665.900 51.400 ;
        RECT 615.600 50.800 665.900 51.000 ;
        RECT 834.100 51.000 884.100 51.400 ;
        RECT 834.100 50.800 884.400 51.000 ;
        RECT 615.600 50.400 665.600 50.800 ;
        RECT 615.400 50.200 665.600 50.400 ;
        RECT 834.400 50.400 884.400 50.800 ;
        RECT 834.400 50.200 884.600 50.400 ;
        RECT 615.400 49.800 665.400 50.200 ;
        RECT 615.200 49.600 665.400 49.800 ;
        RECT 834.600 49.800 884.600 50.200 ;
        RECT 834.600 49.600 884.800 49.800 ;
        RECT 615.200 49.200 665.200 49.600 ;
        RECT 615.000 49.000 665.200 49.200 ;
        RECT 834.800 49.200 884.800 49.600 ;
        RECT 834.800 49.000 885.000 49.200 ;
        RECT 615.000 48.600 665.000 49.000 ;
        RECT 614.800 48.400 665.000 48.600 ;
        RECT 835.000 48.600 885.000 49.000 ;
        RECT 835.000 48.400 885.200 48.600 ;
        RECT 614.800 48.000 664.800 48.400 ;
        RECT 614.500 47.800 664.800 48.000 ;
        RECT 835.200 48.000 885.200 48.400 ;
        RECT 835.200 47.800 885.500 48.000 ;
        RECT 614.500 47.400 664.500 47.800 ;
        RECT 614.300 47.200 664.500 47.400 ;
        RECT 835.500 47.400 885.500 47.800 ;
        RECT 835.500 47.200 885.700 47.400 ;
        RECT 614.300 46.800 664.300 47.200 ;
        RECT 614.100 46.600 664.300 46.800 ;
        RECT 835.700 46.800 885.700 47.200 ;
        RECT 835.700 46.600 885.900 46.800 ;
        RECT 614.100 46.200 664.100 46.600 ;
        RECT 613.800 46.000 664.100 46.200 ;
        RECT 835.900 46.200 885.900 46.600 ;
        RECT 835.900 46.000 886.200 46.200 ;
        RECT 613.800 45.600 663.800 46.000 ;
        RECT 613.600 45.400 663.800 45.600 ;
        RECT 836.200 45.600 886.200 46.000 ;
        RECT 836.200 45.400 886.400 45.600 ;
        RECT 613.600 45.000 663.600 45.400 ;
        RECT 613.400 44.800 663.600 45.000 ;
        RECT 836.400 45.000 886.400 45.400 ;
        RECT 836.400 44.800 886.600 45.000 ;
        RECT 613.400 44.400 663.400 44.800 ;
        RECT 613.200 44.200 663.400 44.400 ;
        RECT 836.600 44.400 886.600 44.800 ;
        RECT 836.600 44.200 886.800 44.400 ;
        RECT 613.200 43.800 663.200 44.200 ;
        RECT 613.000 43.600 663.200 43.800 ;
        RECT 836.800 43.800 886.800 44.200 ;
        RECT 836.800 43.600 887.000 43.800 ;
        RECT 613.000 43.200 663.000 43.600 ;
        RECT 612.700 43.000 663.000 43.200 ;
        RECT 837.000 43.200 887.000 43.600 ;
        RECT 837.000 43.000 887.300 43.200 ;
        RECT 612.700 42.600 662.700 43.000 ;
        RECT 612.500 42.400 662.700 42.600 ;
        RECT 837.300 42.600 887.300 43.000 ;
        RECT 837.300 42.400 887.500 42.600 ;
        RECT 612.500 42.000 662.500 42.400 ;
        RECT 612.300 41.800 662.500 42.000 ;
        RECT 837.500 42.000 887.500 42.400 ;
        RECT 837.500 41.800 887.700 42.000 ;
        RECT 612.300 41.400 662.300 41.800 ;
        RECT 612.000 41.200 662.300 41.400 ;
        RECT 837.700 41.400 887.700 41.800 ;
        RECT 837.700 41.200 888.000 41.400 ;
        RECT 612.000 40.800 662.000 41.200 ;
        RECT 611.800 40.600 662.000 40.800 ;
        RECT 838.000 40.800 888.000 41.200 ;
        RECT 838.000 40.600 888.200 40.800 ;
        RECT 611.800 40.200 661.800 40.600 ;
        RECT 611.600 40.000 661.800 40.200 ;
        RECT 838.200 40.200 888.200 40.600 ;
        RECT 838.200 40.000 888.400 40.200 ;
        RECT 611.600 39.600 661.600 40.000 ;
        RECT 611.400 39.400 661.600 39.600 ;
        RECT 838.400 39.600 888.400 40.000 ;
        RECT 838.400 39.400 888.600 39.600 ;
        RECT 611.400 39.000 661.400 39.400 ;
        RECT 611.200 38.800 661.400 39.000 ;
        RECT 838.600 39.000 888.600 39.400 ;
        RECT 838.600 38.800 888.800 39.000 ;
        RECT 611.200 38.400 661.200 38.800 ;
        RECT 610.900 38.200 661.200 38.400 ;
        RECT 838.800 38.400 888.800 38.800 ;
        RECT 838.800 38.200 889.100 38.400 ;
        RECT 610.900 37.800 660.900 38.200 ;
        RECT 610.700 37.600 660.900 37.800 ;
        RECT 839.100 37.800 889.100 38.200 ;
        RECT 839.100 37.600 889.300 37.800 ;
        RECT 610.700 37.200 660.700 37.600 ;
        RECT 610.500 37.000 660.700 37.200 ;
        RECT 839.300 37.200 889.300 37.600 ;
        RECT 839.300 37.000 889.500 37.200 ;
        RECT 610.500 36.600 660.500 37.000 ;
        RECT 610.200 36.400 660.500 36.600 ;
        RECT 839.500 36.600 889.500 37.000 ;
        RECT 839.500 36.400 889.800 36.600 ;
        RECT 610.200 36.000 660.200 36.400 ;
        RECT 610.000 35.800 660.200 36.000 ;
        RECT 839.800 36.000 889.800 36.400 ;
        RECT 839.800 35.800 890.000 36.000 ;
        RECT 610.000 35.400 660.000 35.800 ;
        RECT 609.800 35.200 660.000 35.400 ;
        RECT 840.000 35.400 890.000 35.800 ;
        RECT 840.000 35.200 890.200 35.400 ;
        RECT 609.800 34.800 659.800 35.200 ;
        RECT 609.600 34.600 659.800 34.800 ;
        RECT 840.200 34.800 890.200 35.200 ;
        RECT 840.200 34.600 890.400 34.800 ;
        RECT 609.600 34.200 659.600 34.600 ;
        RECT 609.400 34.000 659.600 34.200 ;
        RECT 840.400 34.200 890.400 34.600 ;
        RECT 840.400 34.000 890.600 34.200 ;
        RECT 609.400 33.600 659.400 34.000 ;
        RECT 609.100 33.400 659.400 33.600 ;
        RECT 840.600 33.600 890.600 34.000 ;
        RECT 840.600 33.400 890.900 33.600 ;
        RECT 609.100 33.000 659.100 33.400 ;
        RECT 608.900 32.800 659.100 33.000 ;
        RECT 840.900 33.000 890.900 33.400 ;
        RECT 840.900 32.800 891.100 33.000 ;
        RECT 608.900 32.400 658.900 32.800 ;
        RECT 608.700 32.200 658.900 32.400 ;
        RECT 841.100 32.400 891.100 32.800 ;
        RECT 841.100 32.200 891.300 32.400 ;
        RECT 608.700 31.800 658.700 32.200 ;
        RECT 608.400 31.600 658.700 31.800 ;
        RECT 841.300 31.800 891.300 32.200 ;
        RECT 841.300 31.600 891.600 31.800 ;
        RECT 608.400 31.200 658.400 31.600 ;
        RECT 608.200 31.000 658.400 31.200 ;
        RECT 841.600 31.200 891.600 31.600 ;
        RECT 841.600 31.000 891.800 31.200 ;
        RECT 608.200 30.600 658.200 31.000 ;
        RECT 608.000 30.400 658.200 30.600 ;
        RECT 841.800 30.600 891.800 31.000 ;
        RECT 841.800 30.400 892.000 30.600 ;
        RECT 608.000 30.000 658.000 30.400 ;
        RECT 607.800 29.800 658.000 30.000 ;
        RECT 842.000 30.000 892.000 30.400 ;
        RECT 842.000 29.800 892.200 30.000 ;
        RECT 607.800 29.400 657.800 29.800 ;
        RECT 607.600 29.200 657.800 29.400 ;
        RECT 842.200 29.400 892.200 29.800 ;
        RECT 842.200 29.200 892.400 29.400 ;
        RECT 607.600 28.800 657.600 29.200 ;
        RECT 607.300 28.600 657.600 28.800 ;
        RECT 842.400 28.800 892.400 29.200 ;
        RECT 842.400 28.600 892.700 28.800 ;
        RECT 607.300 28.200 657.300 28.600 ;
        RECT 607.100 28.000 657.300 28.200 ;
        RECT 842.700 28.200 892.700 28.600 ;
        RECT 842.700 28.000 892.900 28.200 ;
        RECT 607.100 27.600 657.100 28.000 ;
        RECT 606.900 27.400 657.100 27.600 ;
        RECT 842.900 27.600 892.900 28.000 ;
        RECT 842.900 27.400 893.100 27.600 ;
        RECT 606.900 27.000 656.900 27.400 ;
        RECT 606.600 26.800 656.900 27.000 ;
        RECT 843.100 27.000 893.100 27.400 ;
        RECT 843.100 26.800 893.400 27.000 ;
        RECT 606.600 26.400 656.600 26.800 ;
        RECT 606.400 26.200 656.600 26.400 ;
        RECT 843.400 26.400 893.400 26.800 ;
        RECT 843.400 26.200 893.600 26.400 ;
        RECT 606.400 25.800 656.400 26.200 ;
        RECT 606.200 25.600 656.400 25.800 ;
        RECT 843.600 25.800 893.600 26.200 ;
        RECT 843.600 25.600 893.800 25.800 ;
        RECT 606.200 25.200 656.200 25.600 ;
        RECT 606.000 25.000 656.200 25.200 ;
        RECT 843.800 25.200 893.800 25.600 ;
        RECT 843.800 25.000 894.000 25.200 ;
        RECT 606.000 24.600 656.000 25.000 ;
        RECT 605.800 24.400 656.000 24.600 ;
        RECT 844.000 24.600 894.000 25.000 ;
        RECT 844.000 24.400 894.200 24.600 ;
        RECT 605.800 24.000 655.800 24.400 ;
        RECT 605.500 23.800 655.800 24.000 ;
        RECT 844.200 24.000 894.200 24.400 ;
        RECT 844.200 23.800 894.500 24.000 ;
        RECT 605.500 23.400 655.500 23.800 ;
        RECT 605.300 23.200 655.500 23.400 ;
        RECT 844.500 23.400 894.500 23.800 ;
        RECT 844.500 23.200 894.700 23.400 ;
        RECT 605.300 22.800 655.300 23.200 ;
        RECT 605.100 22.600 655.300 22.800 ;
        RECT 844.700 22.800 894.700 23.200 ;
        RECT 844.700 22.600 894.900 22.800 ;
        RECT 605.100 22.200 655.100 22.600 ;
        RECT 604.800 22.000 655.100 22.200 ;
        RECT 844.900 22.200 894.900 22.600 ;
        RECT 844.900 22.000 895.200 22.200 ;
        RECT 604.800 21.600 654.800 22.000 ;
        RECT 604.600 21.400 654.800 21.600 ;
        RECT 845.200 21.600 895.200 22.000 ;
        RECT 845.200 21.400 895.400 21.600 ;
        RECT 604.600 21.000 654.600 21.400 ;
        RECT 604.400 20.800 654.600 21.000 ;
        RECT 845.400 21.000 895.400 21.400 ;
        RECT 845.400 20.800 895.600 21.000 ;
        RECT 604.400 20.400 654.400 20.800 ;
        RECT 604.200 20.200 654.400 20.400 ;
        RECT 845.600 20.400 895.600 20.800 ;
        RECT 845.600 20.200 895.800 20.400 ;
        RECT 604.200 19.800 654.200 20.200 ;
        RECT 604.000 19.600 654.200 19.800 ;
        RECT 845.800 19.800 895.800 20.200 ;
        RECT 845.800 19.600 896.000 19.800 ;
        RECT 604.000 19.200 654.000 19.600 ;
        RECT 603.700 19.000 654.000 19.200 ;
        RECT 846.000 19.200 896.000 19.600 ;
        RECT 846.000 19.000 896.300 19.200 ;
        RECT 603.700 18.600 653.700 19.000 ;
        RECT 603.500 18.400 653.700 18.600 ;
        RECT 846.300 18.600 896.300 19.000 ;
        RECT 846.300 18.400 896.500 18.600 ;
        RECT 603.500 18.000 653.500 18.400 ;
        RECT 603.300 17.800 653.500 18.000 ;
        RECT 846.500 18.000 896.500 18.400 ;
        RECT 846.500 17.800 896.700 18.000 ;
        RECT 603.300 17.400 653.300 17.800 ;
        RECT 603.000 17.200 653.300 17.400 ;
        RECT 846.700 17.400 896.700 17.800 ;
        RECT 846.700 17.200 897.000 17.400 ;
        RECT 603.000 16.800 653.000 17.200 ;
        RECT 602.800 16.600 653.000 16.800 ;
        RECT 847.000 16.800 897.000 17.200 ;
        RECT 847.000 16.600 897.200 16.800 ;
        RECT 602.800 16.200 652.800 16.600 ;
        RECT 602.600 16.000 652.800 16.200 ;
        RECT 847.200 16.200 897.200 16.600 ;
        RECT 847.200 16.000 897.400 16.200 ;
        RECT 602.600 15.600 652.600 16.000 ;
        RECT 602.400 15.400 652.600 15.600 ;
        RECT 847.400 15.600 897.400 16.000 ;
        RECT 847.400 15.400 897.600 15.600 ;
        RECT 602.400 15.000 652.400 15.400 ;
        RECT 602.200 14.800 652.400 15.000 ;
        RECT 847.600 15.000 897.600 15.400 ;
        RECT 847.600 14.800 897.800 15.000 ;
        RECT 602.200 14.400 652.200 14.800 ;
        RECT 601.900 14.200 652.200 14.400 ;
        RECT 847.800 14.400 897.800 14.800 ;
        RECT 847.800 14.200 898.100 14.400 ;
        RECT 601.900 13.800 651.900 14.200 ;
        RECT 601.700 13.600 651.900 13.800 ;
        RECT 848.100 13.800 898.100 14.200 ;
        RECT 848.100 13.600 898.300 13.800 ;
        RECT 601.700 13.200 651.700 13.600 ;
        RECT 601.500 13.000 651.700 13.200 ;
        RECT 848.300 13.200 898.300 13.600 ;
        RECT 848.300 13.000 898.500 13.200 ;
        RECT 601.500 12.400 651.500 13.000 ;
        RECT 848.500 12.400 898.500 13.000 ;
        RECT 915.000 12.400 965.000 266.800 ;
        RECT 965.400 266.400 1015.400 266.800 ;
        RECT 965.400 266.200 1015.800 266.400 ;
        RECT 965.800 265.800 1015.800 266.200 ;
        RECT 965.800 265.600 1016.200 265.800 ;
        RECT 966.200 265.200 1016.200 265.600 ;
        RECT 966.200 265.000 1016.600 265.200 ;
        RECT 966.600 264.600 1016.600 265.000 ;
        RECT 966.600 264.400 1017.000 264.600 ;
        RECT 967.000 264.000 1017.000 264.400 ;
        RECT 967.000 263.800 1017.400 264.000 ;
        RECT 967.400 263.400 1017.400 263.800 ;
        RECT 967.400 263.200 1017.800 263.400 ;
        RECT 967.800 262.800 1017.800 263.200 ;
        RECT 967.800 262.600 1018.200 262.800 ;
        RECT 968.200 262.200 1018.200 262.600 ;
        RECT 968.200 262.000 1018.600 262.200 ;
        RECT 968.600 261.600 1018.600 262.000 ;
        RECT 968.600 261.400 1019.000 261.600 ;
        RECT 969.000 261.000 1019.000 261.400 ;
        RECT 969.000 260.800 1019.400 261.000 ;
        RECT 969.400 260.400 1019.400 260.800 ;
        RECT 969.400 260.200 1019.800 260.400 ;
        RECT 969.800 259.800 1019.800 260.200 ;
        RECT 969.800 259.600 1020.200 259.800 ;
        RECT 970.200 259.200 1020.200 259.600 ;
        RECT 970.200 259.000 1020.600 259.200 ;
        RECT 970.600 258.600 1020.600 259.000 ;
        RECT 970.600 258.400 1021.000 258.600 ;
        RECT 971.000 258.000 1021.000 258.400 ;
        RECT 971.000 257.800 1021.400 258.000 ;
        RECT 971.400 257.400 1021.400 257.800 ;
        RECT 971.400 257.200 1021.800 257.400 ;
        RECT 971.800 256.800 1021.800 257.200 ;
        RECT 971.800 256.600 1022.200 256.800 ;
        RECT 972.200 256.200 1022.200 256.600 ;
        RECT 972.200 256.000 1022.600 256.200 ;
        RECT 972.600 255.600 1022.600 256.000 ;
        RECT 972.600 255.400 1023.000 255.600 ;
        RECT 973.000 255.000 1023.000 255.400 ;
        RECT 973.000 254.800 1023.400 255.000 ;
        RECT 973.400 254.400 1023.400 254.800 ;
        RECT 973.400 254.200 1023.800 254.400 ;
        RECT 973.800 253.800 1023.800 254.200 ;
        RECT 973.800 253.600 1024.200 253.800 ;
        RECT 974.200 253.200 1024.200 253.600 ;
        RECT 974.200 253.000 1024.600 253.200 ;
        RECT 974.600 252.600 1024.600 253.000 ;
        RECT 974.600 252.400 1025.000 252.600 ;
        RECT 975.000 252.000 1025.000 252.400 ;
        RECT 975.000 251.800 1025.400 252.000 ;
        RECT 975.400 251.400 1025.400 251.800 ;
        RECT 975.400 251.200 1025.800 251.400 ;
        RECT 975.800 250.800 1025.800 251.200 ;
        RECT 975.800 250.600 1026.200 250.800 ;
        RECT 976.200 250.200 1026.200 250.600 ;
        RECT 976.200 250.000 1026.600 250.200 ;
        RECT 976.600 249.600 1026.600 250.000 ;
        RECT 976.600 249.400 1027.000 249.600 ;
        RECT 977.000 249.000 1027.000 249.400 ;
        RECT 977.000 248.800 1027.400 249.000 ;
        RECT 977.400 248.400 1027.400 248.800 ;
        RECT 977.400 248.200 1027.800 248.400 ;
        RECT 977.800 247.800 1027.800 248.200 ;
        RECT 977.800 247.600 1028.200 247.800 ;
        RECT 978.200 247.200 1028.200 247.600 ;
        RECT 978.200 247.000 1028.600 247.200 ;
        RECT 978.600 246.600 1028.600 247.000 ;
        RECT 978.600 246.400 1029.000 246.600 ;
        RECT 979.000 246.000 1029.000 246.400 ;
        RECT 979.000 245.800 1029.400 246.000 ;
        RECT 979.400 245.400 1029.400 245.800 ;
        RECT 979.400 245.200 1029.800 245.400 ;
        RECT 979.800 244.800 1029.800 245.200 ;
        RECT 979.800 244.600 1030.200 244.800 ;
        RECT 980.200 244.200 1030.200 244.600 ;
        RECT 980.200 244.000 1030.600 244.200 ;
        RECT 980.600 243.600 1030.600 244.000 ;
        RECT 980.600 243.400 1031.000 243.600 ;
        RECT 981.000 243.000 1031.000 243.400 ;
        RECT 981.000 242.800 1031.400 243.000 ;
        RECT 981.400 242.400 1031.400 242.800 ;
        RECT 981.400 242.200 1031.800 242.400 ;
        RECT 981.800 241.800 1031.800 242.200 ;
        RECT 981.800 241.600 1032.200 241.800 ;
        RECT 982.200 241.200 1032.200 241.600 ;
        RECT 982.200 241.000 1032.600 241.200 ;
        RECT 982.600 240.600 1032.600 241.000 ;
        RECT 982.600 240.400 1033.000 240.600 ;
        RECT 983.000 240.000 1033.000 240.400 ;
        RECT 983.000 239.800 1033.400 240.000 ;
        RECT 983.400 239.400 1033.400 239.800 ;
        RECT 983.400 239.200 1033.800 239.400 ;
        RECT 983.800 238.800 1033.800 239.200 ;
        RECT 983.800 238.600 1034.200 238.800 ;
        RECT 984.200 238.200 1034.200 238.600 ;
        RECT 984.200 238.000 1034.600 238.200 ;
        RECT 984.600 237.600 1034.600 238.000 ;
        RECT 984.600 237.400 1035.000 237.600 ;
        RECT 985.000 237.000 1035.000 237.400 ;
        RECT 985.000 236.800 1035.400 237.000 ;
        RECT 985.400 236.400 1035.400 236.800 ;
        RECT 985.400 236.200 1035.800 236.400 ;
        RECT 985.800 235.800 1035.800 236.200 ;
        RECT 985.800 235.600 1036.200 235.800 ;
        RECT 986.200 235.200 1036.200 235.600 ;
        RECT 986.200 235.000 1036.600 235.200 ;
        RECT 986.600 234.600 1036.600 235.000 ;
        RECT 986.600 234.400 1037.000 234.600 ;
        RECT 987.000 234.000 1037.000 234.400 ;
        RECT 987.000 233.800 1037.400 234.000 ;
        RECT 987.400 233.400 1037.400 233.800 ;
        RECT 987.400 233.200 1037.800 233.400 ;
        RECT 987.800 232.800 1037.800 233.200 ;
        RECT 987.800 232.600 1038.200 232.800 ;
        RECT 988.200 232.200 1038.200 232.600 ;
        RECT 988.200 232.000 1038.600 232.200 ;
        RECT 988.600 231.600 1038.600 232.000 ;
        RECT 988.600 231.400 1039.000 231.600 ;
        RECT 989.000 231.000 1039.000 231.400 ;
        RECT 989.000 230.800 1039.400 231.000 ;
        RECT 989.400 230.400 1039.400 230.800 ;
        RECT 989.400 230.200 1039.800 230.400 ;
        RECT 989.800 229.800 1039.800 230.200 ;
        RECT 989.800 229.600 1040.200 229.800 ;
        RECT 990.200 229.200 1040.200 229.600 ;
        RECT 990.200 229.000 1040.600 229.200 ;
        RECT 990.600 228.600 1040.600 229.000 ;
        RECT 990.600 228.400 1041.000 228.600 ;
        RECT 991.000 228.000 1041.000 228.400 ;
        RECT 991.000 227.800 1041.400 228.000 ;
        RECT 991.400 227.400 1041.400 227.800 ;
        RECT 991.400 227.200 1041.800 227.400 ;
        RECT 991.800 226.800 1041.800 227.200 ;
        RECT 991.800 226.600 1042.200 226.800 ;
        RECT 992.200 226.200 1042.200 226.600 ;
        RECT 992.200 226.000 1042.600 226.200 ;
        RECT 992.600 225.600 1042.600 226.000 ;
        RECT 992.600 225.400 1043.000 225.600 ;
        RECT 993.000 225.000 1043.000 225.400 ;
        RECT 993.000 224.800 1043.400 225.000 ;
        RECT 993.400 224.400 1043.400 224.800 ;
        RECT 993.400 224.200 1043.800 224.400 ;
        RECT 993.800 223.800 1043.800 224.200 ;
        RECT 993.800 223.600 1044.200 223.800 ;
        RECT 994.200 223.200 1044.200 223.600 ;
        RECT 994.200 223.000 1044.600 223.200 ;
        RECT 994.600 222.600 1044.600 223.000 ;
        RECT 994.600 222.400 1045.000 222.600 ;
        RECT 995.000 222.000 1045.000 222.400 ;
        RECT 995.000 221.800 1045.400 222.000 ;
        RECT 995.400 221.400 1045.400 221.800 ;
        RECT 995.400 221.200 1045.800 221.400 ;
        RECT 995.800 220.800 1045.800 221.200 ;
        RECT 995.800 220.600 1046.200 220.800 ;
        RECT 996.200 220.200 1046.200 220.600 ;
        RECT 996.200 220.000 1046.600 220.200 ;
        RECT 996.600 219.600 1046.600 220.000 ;
        RECT 996.600 219.400 1047.000 219.600 ;
        RECT 997.000 219.000 1047.000 219.400 ;
        RECT 997.000 218.800 1047.400 219.000 ;
        RECT 997.400 218.400 1047.400 218.800 ;
        RECT 997.400 218.200 1047.800 218.400 ;
        RECT 997.800 217.800 1047.800 218.200 ;
        RECT 997.800 217.600 1048.200 217.800 ;
        RECT 998.200 217.200 1048.200 217.600 ;
        RECT 998.200 217.000 1048.600 217.200 ;
        RECT 998.600 216.600 1048.600 217.000 ;
        RECT 998.600 216.400 1049.000 216.600 ;
        RECT 999.000 216.000 1049.000 216.400 ;
        RECT 999.000 215.800 1049.400 216.000 ;
        RECT 999.400 215.400 1049.400 215.800 ;
        RECT 999.400 215.200 1049.800 215.400 ;
        RECT 999.800 214.800 1049.800 215.200 ;
        RECT 999.800 214.600 1050.200 214.800 ;
        RECT 1000.200 214.200 1050.200 214.600 ;
        RECT 1000.200 214.000 1050.600 214.200 ;
        RECT 1000.600 213.600 1050.600 214.000 ;
        RECT 1000.600 213.400 1051.000 213.600 ;
        RECT 1001.000 213.000 1051.000 213.400 ;
        RECT 1001.000 212.800 1051.400 213.000 ;
        RECT 1001.400 212.400 1051.400 212.800 ;
        RECT 1001.400 212.200 1051.800 212.400 ;
        RECT 1001.800 211.800 1051.800 212.200 ;
        RECT 1001.800 211.600 1052.200 211.800 ;
        RECT 1002.200 211.200 1052.200 211.600 ;
        RECT 1002.200 211.000 1052.600 211.200 ;
        RECT 1002.600 210.600 1052.600 211.000 ;
        RECT 1002.600 210.400 1053.000 210.600 ;
        RECT 1003.000 210.000 1053.000 210.400 ;
        RECT 1003.000 209.800 1053.400 210.000 ;
        RECT 1003.400 209.400 1053.400 209.800 ;
        RECT 1003.400 209.200 1053.800 209.400 ;
        RECT 1003.800 208.800 1053.800 209.200 ;
        RECT 1003.800 208.600 1054.200 208.800 ;
        RECT 1004.200 208.200 1054.200 208.600 ;
        RECT 1004.200 208.000 1054.600 208.200 ;
        RECT 1004.600 207.600 1054.600 208.000 ;
        RECT 1004.600 207.400 1055.000 207.600 ;
        RECT 1005.000 207.000 1055.000 207.400 ;
        RECT 1005.000 206.800 1055.400 207.000 ;
        RECT 1005.400 206.400 1055.400 206.800 ;
        RECT 1005.400 206.200 1055.800 206.400 ;
        RECT 1005.800 205.800 1055.800 206.200 ;
        RECT 1005.800 205.600 1056.200 205.800 ;
        RECT 1006.200 205.200 1056.200 205.600 ;
        RECT 1006.200 205.000 1056.600 205.200 ;
        RECT 1006.600 204.600 1056.600 205.000 ;
        RECT 1006.600 204.400 1057.000 204.600 ;
        RECT 1007.000 204.000 1057.000 204.400 ;
        RECT 1007.000 203.800 1057.400 204.000 ;
        RECT 1007.400 203.400 1057.400 203.800 ;
        RECT 1007.400 203.200 1057.800 203.400 ;
        RECT 1007.800 202.800 1057.800 203.200 ;
        RECT 1007.800 202.600 1058.200 202.800 ;
        RECT 1008.200 202.200 1058.200 202.600 ;
        RECT 1008.200 202.000 1058.600 202.200 ;
        RECT 1008.600 201.600 1058.600 202.000 ;
        RECT 1008.600 201.400 1059.000 201.600 ;
        RECT 1009.000 201.000 1059.000 201.400 ;
        RECT 1009.000 200.800 1059.400 201.000 ;
        RECT 1009.400 200.400 1059.400 200.800 ;
        RECT 1009.400 200.200 1059.800 200.400 ;
        RECT 1009.800 199.800 1059.800 200.200 ;
        RECT 1009.800 199.600 1060.200 199.800 ;
        RECT 1010.200 199.200 1060.200 199.600 ;
        RECT 1010.200 199.000 1060.600 199.200 ;
        RECT 1010.600 198.600 1060.600 199.000 ;
        RECT 1010.600 198.400 1061.000 198.600 ;
        RECT 1011.000 198.000 1061.000 198.400 ;
        RECT 1011.000 197.800 1061.400 198.000 ;
        RECT 1011.400 197.400 1061.400 197.800 ;
        RECT 1011.400 197.200 1061.800 197.400 ;
        RECT 1011.800 196.800 1061.800 197.200 ;
        RECT 1011.800 196.600 1062.200 196.800 ;
        RECT 1012.200 196.200 1062.200 196.600 ;
        RECT 1012.200 196.000 1062.600 196.200 ;
        RECT 1012.600 195.600 1062.600 196.000 ;
        RECT 1012.600 195.400 1063.000 195.600 ;
        RECT 1013.000 195.000 1063.000 195.400 ;
        RECT 1013.000 194.800 1063.400 195.000 ;
        RECT 1013.400 194.400 1063.400 194.800 ;
        RECT 1013.400 194.200 1063.800 194.400 ;
        RECT 1013.800 193.800 1063.800 194.200 ;
        RECT 1013.800 193.600 1064.200 193.800 ;
        RECT 1014.200 193.200 1064.200 193.600 ;
        RECT 1014.200 193.000 1064.600 193.200 ;
        RECT 1014.600 192.600 1064.600 193.000 ;
        RECT 1014.600 192.400 1065.000 192.600 ;
        RECT 1015.000 192.000 1065.000 192.400 ;
        RECT 1015.000 191.800 1065.400 192.000 ;
        RECT 1015.400 191.400 1065.400 191.800 ;
        RECT 1015.400 191.200 1065.800 191.400 ;
        RECT 1015.800 190.800 1065.800 191.200 ;
        RECT 1015.800 190.600 1066.200 190.800 ;
        RECT 1016.200 190.200 1066.200 190.600 ;
        RECT 1016.200 190.000 1066.600 190.200 ;
        RECT 1016.600 189.600 1066.600 190.000 ;
        RECT 1016.600 189.400 1067.000 189.600 ;
        RECT 1017.000 189.000 1067.000 189.400 ;
        RECT 1017.000 188.800 1067.400 189.000 ;
        RECT 1017.400 188.400 1067.400 188.800 ;
        RECT 1017.400 188.200 1067.800 188.400 ;
        RECT 1017.800 187.800 1067.800 188.200 ;
        RECT 1017.800 187.600 1068.200 187.800 ;
        RECT 1018.200 187.200 1068.200 187.600 ;
        RECT 1018.200 187.000 1068.600 187.200 ;
        RECT 1018.600 186.600 1068.600 187.000 ;
        RECT 1018.600 186.400 1069.000 186.600 ;
        RECT 1019.000 186.000 1069.000 186.400 ;
        RECT 1019.000 185.800 1069.400 186.000 ;
        RECT 1019.400 185.400 1069.400 185.800 ;
        RECT 1019.400 185.200 1069.800 185.400 ;
        RECT 1019.800 184.800 1069.800 185.200 ;
        RECT 1019.800 184.600 1070.200 184.800 ;
        RECT 1020.200 184.200 1070.200 184.600 ;
        RECT 1020.200 184.000 1070.600 184.200 ;
        RECT 1020.600 183.600 1070.600 184.000 ;
        RECT 1020.600 183.400 1071.000 183.600 ;
        RECT 1021.000 183.000 1071.000 183.400 ;
        RECT 1021.000 182.800 1071.400 183.000 ;
        RECT 1021.400 182.400 1071.400 182.800 ;
        RECT 1021.400 182.200 1071.800 182.400 ;
        RECT 1021.800 181.800 1071.800 182.200 ;
        RECT 1021.800 181.600 1072.200 181.800 ;
        RECT 1022.200 181.200 1072.200 181.600 ;
        RECT 1022.200 181.000 1072.600 181.200 ;
        RECT 1022.600 180.600 1072.600 181.000 ;
        RECT 1022.600 180.400 1073.000 180.600 ;
        RECT 1023.000 180.000 1073.000 180.400 ;
        RECT 1023.000 179.800 1073.400 180.000 ;
        RECT 1023.400 179.400 1073.400 179.800 ;
        RECT 1023.400 179.200 1073.800 179.400 ;
        RECT 1023.800 178.800 1073.800 179.200 ;
        RECT 1023.800 178.600 1074.200 178.800 ;
        RECT 1024.200 178.200 1074.200 178.600 ;
        RECT 1024.200 178.000 1074.600 178.200 ;
        RECT 1024.600 177.600 1074.600 178.000 ;
        RECT 1024.600 177.400 1075.000 177.600 ;
        RECT 1025.000 177.000 1075.000 177.400 ;
        RECT 1025.000 176.800 1075.400 177.000 ;
        RECT 1025.400 176.400 1075.400 176.800 ;
        RECT 1025.400 176.200 1075.800 176.400 ;
        RECT 1025.800 175.800 1075.800 176.200 ;
        RECT 1025.800 175.600 1076.200 175.800 ;
        RECT 1026.200 175.200 1076.200 175.600 ;
        RECT 1026.200 175.000 1076.600 175.200 ;
        RECT 1026.600 174.600 1076.600 175.000 ;
        RECT 1026.600 174.400 1077.000 174.600 ;
        RECT 1027.000 174.000 1077.000 174.400 ;
        RECT 1027.000 173.800 1077.400 174.000 ;
        RECT 1027.400 173.400 1077.400 173.800 ;
        RECT 1027.400 173.200 1077.800 173.400 ;
        RECT 1027.800 172.800 1077.800 173.200 ;
        RECT 1027.800 172.600 1078.200 172.800 ;
        RECT 1028.200 172.200 1078.200 172.600 ;
        RECT 1028.200 172.000 1078.600 172.200 ;
        RECT 1028.600 171.600 1078.600 172.000 ;
        RECT 1028.600 171.400 1079.000 171.600 ;
        RECT 1029.000 171.000 1079.000 171.400 ;
        RECT 1029.000 170.800 1079.400 171.000 ;
        RECT 1029.400 170.400 1079.400 170.800 ;
        RECT 1029.400 170.200 1079.800 170.400 ;
        RECT 1029.800 169.800 1079.800 170.200 ;
        RECT 1029.800 169.600 1080.200 169.800 ;
        RECT 1030.200 169.200 1080.200 169.600 ;
        RECT 1030.200 169.000 1080.600 169.200 ;
        RECT 1030.600 168.600 1080.600 169.000 ;
        RECT 1030.600 168.400 1081.000 168.600 ;
        RECT 1031.000 168.000 1081.000 168.400 ;
        RECT 1031.000 167.800 1081.400 168.000 ;
        RECT 1031.400 167.400 1081.400 167.800 ;
        RECT 1031.400 167.200 1081.800 167.400 ;
        RECT 1031.800 166.800 1081.800 167.200 ;
        RECT 1031.800 166.600 1082.200 166.800 ;
        RECT 1032.200 166.200 1082.200 166.600 ;
        RECT 1032.200 166.000 1082.600 166.200 ;
        RECT 1032.600 165.600 1082.600 166.000 ;
        RECT 1032.600 165.400 1083.000 165.600 ;
        RECT 1033.000 165.000 1083.000 165.400 ;
        RECT 1033.000 164.800 1083.400 165.000 ;
        RECT 1033.400 164.400 1083.400 164.800 ;
        RECT 1033.400 164.200 1083.800 164.400 ;
        RECT 1033.800 163.800 1083.800 164.200 ;
        RECT 1033.800 163.600 1084.200 163.800 ;
        RECT 1034.200 163.200 1084.200 163.600 ;
        RECT 1034.200 163.000 1084.600 163.200 ;
        RECT 1034.600 162.600 1084.600 163.000 ;
        RECT 1034.600 162.400 1085.000 162.600 ;
        RECT 1035.000 162.000 1085.000 162.400 ;
        RECT 1035.000 161.800 1085.400 162.000 ;
        RECT 1035.400 161.400 1085.400 161.800 ;
        RECT 1035.400 161.200 1085.800 161.400 ;
        RECT 1035.800 160.800 1085.800 161.200 ;
        RECT 1035.800 160.600 1086.200 160.800 ;
        RECT 1036.200 160.200 1086.200 160.600 ;
        RECT 1036.200 160.000 1086.600 160.200 ;
        RECT 1036.600 159.600 1086.600 160.000 ;
        RECT 1036.600 159.400 1087.000 159.600 ;
        RECT 1037.000 159.000 1087.000 159.400 ;
        RECT 1037.000 158.800 1087.400 159.000 ;
        RECT 1037.400 158.400 1087.400 158.800 ;
        RECT 1037.400 158.200 1087.800 158.400 ;
        RECT 1037.800 157.800 1087.800 158.200 ;
        RECT 1037.800 157.600 1088.200 157.800 ;
        RECT 1038.200 157.200 1088.200 157.600 ;
        RECT 1038.200 157.000 1088.600 157.200 ;
        RECT 1038.600 156.600 1088.600 157.000 ;
        RECT 1038.600 156.400 1089.000 156.600 ;
        RECT 1039.000 156.000 1089.000 156.400 ;
        RECT 1039.000 155.800 1089.400 156.000 ;
        RECT 1039.400 155.400 1089.400 155.800 ;
        RECT 1039.400 155.200 1089.800 155.400 ;
        RECT 1039.800 154.800 1089.800 155.200 ;
        RECT 1039.800 154.600 1090.200 154.800 ;
        RECT 1040.200 154.200 1090.200 154.600 ;
        RECT 1040.200 154.000 1090.600 154.200 ;
        RECT 1040.600 153.600 1090.600 154.000 ;
        RECT 1040.600 153.400 1091.000 153.600 ;
        RECT 1041.000 153.000 1091.000 153.400 ;
        RECT 1041.000 152.800 1091.400 153.000 ;
        RECT 1041.400 152.400 1091.400 152.800 ;
        RECT 1041.400 152.200 1091.800 152.400 ;
        RECT 1041.800 151.800 1091.800 152.200 ;
        RECT 1041.800 151.600 1092.200 151.800 ;
        RECT 1042.200 151.200 1092.200 151.600 ;
        RECT 1042.200 151.000 1092.600 151.200 ;
        RECT 1042.600 150.600 1092.600 151.000 ;
        RECT 1042.600 150.400 1093.000 150.600 ;
        RECT 1043.000 150.000 1093.000 150.400 ;
        RECT 1043.000 149.800 1093.400 150.000 ;
        RECT 1043.400 149.400 1093.400 149.800 ;
        RECT 1043.400 149.200 1093.800 149.400 ;
        RECT 1043.800 148.800 1093.800 149.200 ;
        RECT 1043.800 148.600 1094.200 148.800 ;
        RECT 1044.200 148.200 1094.200 148.600 ;
        RECT 1044.200 148.000 1094.600 148.200 ;
        RECT 1044.600 147.600 1094.600 148.000 ;
        RECT 1044.600 147.400 1095.000 147.600 ;
        RECT 1045.000 147.000 1095.000 147.400 ;
        RECT 1045.000 146.800 1095.400 147.000 ;
        RECT 1045.400 146.400 1095.400 146.800 ;
        RECT 1045.400 146.200 1095.800 146.400 ;
        RECT 1045.800 145.800 1095.800 146.200 ;
        RECT 1045.800 145.600 1096.200 145.800 ;
        RECT 1046.200 145.200 1096.200 145.600 ;
        RECT 1046.200 145.000 1096.600 145.200 ;
        RECT 1046.600 144.600 1096.600 145.000 ;
        RECT 1046.600 144.400 1097.000 144.600 ;
        RECT 1047.000 144.000 1097.000 144.400 ;
        RECT 1047.000 143.800 1097.400 144.000 ;
        RECT 1047.400 143.400 1097.400 143.800 ;
        RECT 1047.400 143.200 1097.800 143.400 ;
        RECT 1047.800 142.800 1097.800 143.200 ;
        RECT 1047.800 142.600 1098.200 142.800 ;
        RECT 1048.200 142.200 1098.200 142.600 ;
        RECT 1048.200 142.000 1098.600 142.200 ;
        RECT 1048.600 141.600 1098.600 142.000 ;
        RECT 1048.600 141.400 1099.000 141.600 ;
        RECT 1049.000 141.000 1099.000 141.400 ;
        RECT 1049.000 140.800 1099.400 141.000 ;
        RECT 1049.400 140.400 1099.400 140.800 ;
        RECT 1049.400 140.200 1099.800 140.400 ;
        RECT 1049.800 139.800 1099.800 140.200 ;
        RECT 1049.800 139.600 1100.200 139.800 ;
        RECT 1050.200 139.200 1100.200 139.600 ;
        RECT 1050.200 139.000 1100.600 139.200 ;
        RECT 1050.600 138.600 1100.600 139.000 ;
        RECT 1050.600 138.400 1101.000 138.600 ;
        RECT 1051.000 138.000 1101.000 138.400 ;
        RECT 1051.000 137.800 1101.400 138.000 ;
        RECT 1051.400 137.400 1101.400 137.800 ;
        RECT 1051.400 137.200 1101.800 137.400 ;
        RECT 1051.800 136.800 1101.800 137.200 ;
        RECT 1051.800 136.600 1102.200 136.800 ;
        RECT 1052.200 136.200 1102.200 136.600 ;
        RECT 1052.200 136.000 1102.600 136.200 ;
        RECT 1052.600 135.600 1102.600 136.000 ;
        RECT 1052.600 135.400 1103.000 135.600 ;
        RECT 1053.000 135.000 1103.000 135.400 ;
        RECT 1053.000 134.800 1103.400 135.000 ;
        RECT 1053.400 134.400 1103.400 134.800 ;
        RECT 1053.400 134.200 1103.800 134.400 ;
        RECT 1053.800 133.800 1103.800 134.200 ;
        RECT 1053.800 133.600 1104.200 133.800 ;
        RECT 1054.200 133.200 1104.200 133.600 ;
        RECT 1054.200 133.000 1104.600 133.200 ;
        RECT 1054.600 132.600 1104.600 133.000 ;
        RECT 1054.600 132.400 1105.000 132.600 ;
        RECT 1055.000 132.000 1105.000 132.400 ;
        RECT 1055.000 131.800 1105.400 132.000 ;
        RECT 1055.400 131.400 1105.400 131.800 ;
        RECT 1055.400 131.200 1105.800 131.400 ;
        RECT 1055.800 130.800 1105.800 131.200 ;
        RECT 1055.800 130.600 1106.200 130.800 ;
        RECT 1056.200 130.200 1106.200 130.600 ;
        RECT 1056.200 130.000 1106.600 130.200 ;
        RECT 1056.600 129.600 1106.600 130.000 ;
        RECT 1056.600 129.400 1107.000 129.600 ;
        RECT 1057.000 129.000 1107.000 129.400 ;
        RECT 1057.000 128.800 1107.400 129.000 ;
        RECT 1057.400 128.400 1107.400 128.800 ;
        RECT 1057.400 128.200 1107.800 128.400 ;
        RECT 1057.800 127.800 1107.800 128.200 ;
        RECT 1057.800 127.600 1108.200 127.800 ;
        RECT 1058.200 127.200 1108.200 127.600 ;
        RECT 1058.200 127.000 1108.600 127.200 ;
        RECT 1058.600 126.600 1108.600 127.000 ;
        RECT 1058.600 126.400 1109.000 126.600 ;
        RECT 1059.000 126.000 1109.000 126.400 ;
        RECT 1059.000 125.800 1109.400 126.000 ;
        RECT 1059.400 125.400 1109.400 125.800 ;
        RECT 1059.400 125.200 1109.800 125.400 ;
        RECT 1059.800 124.800 1109.800 125.200 ;
        RECT 1059.800 124.600 1110.200 124.800 ;
        RECT 1060.200 124.200 1110.200 124.600 ;
        RECT 1060.200 124.000 1110.600 124.200 ;
        RECT 1060.600 123.600 1110.600 124.000 ;
        RECT 1060.600 123.400 1111.000 123.600 ;
        RECT 1061.000 123.000 1111.000 123.400 ;
        RECT 1061.000 122.800 1111.400 123.000 ;
        RECT 1061.400 122.400 1111.400 122.800 ;
        RECT 1061.400 122.200 1111.800 122.400 ;
        RECT 1061.800 121.800 1111.800 122.200 ;
        RECT 1061.800 121.600 1112.200 121.800 ;
        RECT 1062.200 121.200 1112.200 121.600 ;
        RECT 1062.200 121.000 1112.600 121.200 ;
        RECT 1062.600 120.600 1112.600 121.000 ;
        RECT 1062.600 120.400 1113.000 120.600 ;
        RECT 1063.000 120.000 1113.000 120.400 ;
        RECT 1063.000 119.800 1113.400 120.000 ;
        RECT 1063.400 119.400 1113.400 119.800 ;
        RECT 1063.400 119.200 1113.800 119.400 ;
        RECT 1063.800 118.800 1113.800 119.200 ;
        RECT 1063.800 118.600 1114.200 118.800 ;
        RECT 1064.200 118.200 1114.200 118.600 ;
        RECT 1064.200 118.000 1114.600 118.200 ;
        RECT 1064.600 117.600 1114.600 118.000 ;
        RECT 1064.600 117.400 1115.000 117.600 ;
        RECT 1065.000 117.000 1115.000 117.400 ;
        RECT 1065.000 116.800 1115.400 117.000 ;
        RECT 1065.400 116.400 1115.400 116.800 ;
        RECT 1065.400 116.200 1115.800 116.400 ;
        RECT 1065.800 115.800 1115.800 116.200 ;
        RECT 1065.800 115.600 1116.200 115.800 ;
        RECT 1066.200 115.200 1116.200 115.600 ;
        RECT 1066.200 115.000 1116.600 115.200 ;
        RECT 1066.600 114.600 1116.600 115.000 ;
        RECT 1066.600 114.400 1117.000 114.600 ;
        RECT 1067.000 114.000 1117.000 114.400 ;
        RECT 1067.000 113.800 1117.400 114.000 ;
        RECT 1067.400 113.400 1117.400 113.800 ;
        RECT 1067.400 113.200 1117.800 113.400 ;
        RECT 1067.800 112.800 1117.800 113.200 ;
        RECT 1067.800 112.600 1118.200 112.800 ;
        RECT 1068.200 112.200 1118.200 112.600 ;
        RECT 1068.200 112.000 1118.600 112.200 ;
        RECT 1068.600 111.600 1118.600 112.000 ;
        RECT 1068.600 111.400 1119.000 111.600 ;
        RECT 1069.000 111.000 1119.000 111.400 ;
        RECT 1069.000 110.800 1119.400 111.000 ;
        RECT 1069.400 110.400 1119.400 110.800 ;
        RECT 1069.400 110.200 1119.800 110.400 ;
        RECT 1069.800 109.800 1119.800 110.200 ;
        RECT 1069.800 109.600 1120.200 109.800 ;
        RECT 1070.200 109.200 1120.200 109.600 ;
        RECT 1070.200 109.000 1120.600 109.200 ;
        RECT 1070.600 108.600 1120.600 109.000 ;
        RECT 1070.600 108.400 1121.000 108.600 ;
        RECT 1071.000 108.000 1121.000 108.400 ;
        RECT 1071.000 107.800 1121.400 108.000 ;
        RECT 1071.400 107.400 1121.400 107.800 ;
        RECT 1071.400 107.200 1121.800 107.400 ;
        RECT 1071.800 106.800 1121.800 107.200 ;
        RECT 1071.800 106.600 1122.200 106.800 ;
        RECT 1072.200 106.200 1122.200 106.600 ;
        RECT 1072.200 106.000 1122.600 106.200 ;
        RECT 1072.600 105.600 1122.600 106.000 ;
        RECT 1072.600 105.400 1123.000 105.600 ;
        RECT 1073.000 105.000 1123.000 105.400 ;
        RECT 1073.000 104.800 1123.400 105.000 ;
        RECT 1073.400 104.400 1123.400 104.800 ;
        RECT 1073.400 104.200 1123.800 104.400 ;
        RECT 1073.800 103.800 1123.800 104.200 ;
        RECT 1073.800 103.600 1124.200 103.800 ;
        RECT 1074.200 103.200 1124.200 103.600 ;
        RECT 1074.200 103.000 1124.600 103.200 ;
        RECT 1074.600 102.600 1124.600 103.000 ;
        RECT 1074.600 102.400 1125.000 102.600 ;
        RECT 1075.000 102.000 1125.000 102.400 ;
        RECT 1075.000 101.800 1125.400 102.000 ;
        RECT 1075.400 101.400 1125.400 101.800 ;
        RECT 1075.400 101.200 1125.800 101.400 ;
        RECT 1075.800 100.800 1125.800 101.200 ;
        RECT 1075.800 100.600 1126.200 100.800 ;
        RECT 1076.200 100.200 1126.200 100.600 ;
        RECT 1076.200 100.000 1126.600 100.200 ;
        RECT 1076.600 99.600 1126.600 100.000 ;
        RECT 1076.600 99.400 1127.000 99.600 ;
        RECT 1077.000 99.000 1127.000 99.400 ;
        RECT 1077.000 98.800 1127.400 99.000 ;
        RECT 1077.400 98.400 1127.400 98.800 ;
        RECT 1077.400 98.200 1127.800 98.400 ;
        RECT 1077.800 97.800 1127.800 98.200 ;
        RECT 1077.800 97.600 1128.200 97.800 ;
        RECT 1078.200 97.200 1128.200 97.600 ;
        RECT 1078.200 97.000 1128.600 97.200 ;
        RECT 1078.600 96.600 1128.600 97.000 ;
        RECT 1078.600 96.400 1129.000 96.600 ;
        RECT 1079.000 96.000 1129.000 96.400 ;
        RECT 1079.000 95.800 1129.400 96.000 ;
        RECT 1079.400 95.400 1129.400 95.800 ;
        RECT 1079.400 95.200 1129.800 95.400 ;
        RECT 1079.800 94.800 1129.800 95.200 ;
        RECT 1079.800 94.600 1130.200 94.800 ;
        RECT 1080.200 94.200 1130.200 94.600 ;
        RECT 1080.200 94.000 1130.600 94.200 ;
        RECT 1080.600 93.600 1130.600 94.000 ;
        RECT 1080.600 93.400 1131.000 93.600 ;
        RECT 1081.000 93.000 1131.000 93.400 ;
        RECT 1081.000 92.800 1131.400 93.000 ;
        RECT 1081.400 92.400 1131.400 92.800 ;
        RECT 1081.400 92.200 1131.800 92.400 ;
        RECT 1081.800 91.800 1131.800 92.200 ;
        RECT 1081.800 91.600 1132.200 91.800 ;
        RECT 1082.200 91.200 1132.200 91.600 ;
        RECT 1082.200 91.000 1132.600 91.200 ;
        RECT 1082.600 90.600 1132.600 91.000 ;
        RECT 1082.600 90.400 1133.000 90.600 ;
        RECT 1083.000 90.000 1133.000 90.400 ;
        RECT 1083.000 89.800 1133.400 90.000 ;
        RECT 1083.400 89.400 1133.400 89.800 ;
        RECT 1083.400 89.200 1133.800 89.400 ;
        RECT 1083.800 88.800 1133.800 89.200 ;
        RECT 1083.800 88.600 1134.200 88.800 ;
        RECT 1084.200 88.200 1134.200 88.600 ;
        RECT 1084.200 88.000 1134.600 88.200 ;
        RECT 1084.600 87.600 1134.600 88.000 ;
        RECT 1135.000 87.600 1185.000 342.600 ;
        RECT 1084.600 87.400 1185.000 87.600 ;
        RECT 1085.000 86.800 1185.000 87.400 ;
        RECT 1085.400 86.200 1185.000 86.800 ;
        RECT 1085.800 85.600 1185.000 86.200 ;
        RECT 1086.200 85.000 1185.000 85.600 ;
        RECT 1086.600 84.400 1185.000 85.000 ;
        RECT 1087.000 83.800 1185.000 84.400 ;
        RECT 1087.400 83.200 1185.000 83.800 ;
        RECT 1087.800 82.600 1185.000 83.200 ;
        RECT 1088.200 82.000 1185.000 82.600 ;
        RECT 1088.600 81.400 1185.000 82.000 ;
        RECT 1089.000 80.800 1185.000 81.400 ;
        RECT 1089.400 80.200 1185.000 80.800 ;
        RECT 1089.800 79.600 1185.000 80.200 ;
        RECT 1090.200 79.000 1185.000 79.600 ;
        RECT 1090.600 78.400 1185.000 79.000 ;
        RECT 1091.000 77.800 1185.000 78.400 ;
        RECT 1091.400 77.200 1185.000 77.800 ;
        RECT 1091.800 76.600 1185.000 77.200 ;
        RECT 1092.200 76.000 1185.000 76.600 ;
        RECT 1092.600 75.400 1185.000 76.000 ;
        RECT 1093.000 74.800 1185.000 75.400 ;
        RECT 1093.400 74.200 1185.000 74.800 ;
        RECT 1093.800 73.600 1185.000 74.200 ;
        RECT 1094.200 73.000 1185.000 73.600 ;
        RECT 1094.600 72.400 1185.000 73.000 ;
        RECT 1095.000 71.800 1185.000 72.400 ;
        RECT 1095.400 71.200 1185.000 71.800 ;
        RECT 1095.800 70.600 1185.000 71.200 ;
        RECT 1096.200 70.000 1185.000 70.600 ;
        RECT 1096.600 69.400 1185.000 70.000 ;
        RECT 1097.000 68.800 1185.000 69.400 ;
        RECT 1097.400 68.200 1185.000 68.800 ;
        RECT 1097.800 67.600 1185.000 68.200 ;
        RECT 1098.200 67.000 1185.000 67.600 ;
        RECT 1098.600 66.400 1185.000 67.000 ;
        RECT 1099.000 65.800 1185.000 66.400 ;
        RECT 1099.400 65.200 1185.000 65.800 ;
        RECT 1099.800 64.600 1185.000 65.200 ;
        RECT 1100.200 64.000 1185.000 64.600 ;
        RECT 1100.600 63.400 1185.000 64.000 ;
        RECT 1101.000 62.800 1185.000 63.400 ;
        RECT 1101.400 62.200 1185.000 62.800 ;
        RECT 1101.800 61.600 1185.000 62.200 ;
        RECT 1102.200 61.000 1185.000 61.600 ;
        RECT 1102.600 60.400 1185.000 61.000 ;
        RECT 1103.000 59.800 1185.000 60.400 ;
        RECT 1103.400 59.200 1185.000 59.800 ;
        RECT 1103.800 58.600 1185.000 59.200 ;
        RECT 1104.200 58.000 1185.000 58.600 ;
        RECT 1104.600 57.400 1185.000 58.000 ;
        RECT 1105.000 56.800 1185.000 57.400 ;
        RECT 1105.400 56.200 1185.000 56.800 ;
        RECT 1105.800 55.600 1185.000 56.200 ;
        RECT 1106.200 55.000 1185.000 55.600 ;
        RECT 1106.600 54.400 1185.000 55.000 ;
        RECT 1107.000 53.800 1185.000 54.400 ;
        RECT 1107.400 53.200 1185.000 53.800 ;
        RECT 1107.800 52.600 1185.000 53.200 ;
        RECT 1108.200 52.000 1185.000 52.600 ;
        RECT 1108.600 51.400 1185.000 52.000 ;
        RECT 1109.000 50.800 1185.000 51.400 ;
        RECT 1109.400 50.200 1185.000 50.800 ;
        RECT 1109.800 49.600 1185.000 50.200 ;
        RECT 1110.200 49.000 1185.000 49.600 ;
        RECT 1110.600 48.400 1185.000 49.000 ;
        RECT 1111.000 47.800 1185.000 48.400 ;
        RECT 1111.400 47.200 1185.000 47.800 ;
        RECT 1111.800 46.600 1185.000 47.200 ;
        RECT 1112.200 46.000 1185.000 46.600 ;
        RECT 1112.600 45.400 1185.000 46.000 ;
        RECT 1113.000 44.800 1185.000 45.400 ;
        RECT 1113.400 44.200 1185.000 44.800 ;
        RECT 1113.800 43.600 1185.000 44.200 ;
        RECT 1114.200 43.000 1185.000 43.600 ;
        RECT 1114.600 42.400 1185.000 43.000 ;
        RECT 1115.000 41.800 1185.000 42.400 ;
        RECT 1115.400 41.200 1185.000 41.800 ;
        RECT 1115.800 40.600 1185.000 41.200 ;
        RECT 1116.200 40.000 1185.000 40.600 ;
        RECT 1116.600 39.400 1185.000 40.000 ;
        RECT 1117.000 38.800 1185.000 39.400 ;
        RECT 1117.400 38.200 1185.000 38.800 ;
        RECT 1117.800 37.600 1185.000 38.200 ;
        RECT 1118.200 37.000 1185.000 37.600 ;
        RECT 1118.600 36.400 1185.000 37.000 ;
        RECT 1119.000 35.800 1185.000 36.400 ;
        RECT 1119.400 35.200 1185.000 35.800 ;
        RECT 1119.800 34.600 1185.000 35.200 ;
        RECT 1120.200 34.000 1185.000 34.600 ;
        RECT 1120.600 33.400 1185.000 34.000 ;
        RECT 1121.000 32.800 1185.000 33.400 ;
        RECT 1121.400 32.200 1185.000 32.800 ;
        RECT 1121.800 31.600 1185.000 32.200 ;
        RECT 1122.200 31.000 1185.000 31.600 ;
        RECT 1122.600 30.400 1185.000 31.000 ;
        RECT 1123.000 29.800 1185.000 30.400 ;
        RECT 1123.400 29.200 1185.000 29.800 ;
        RECT 1123.800 28.600 1185.000 29.200 ;
        RECT 1124.200 28.000 1185.000 28.600 ;
        RECT 1124.600 27.400 1185.000 28.000 ;
        RECT 1125.000 26.800 1185.000 27.400 ;
        RECT 1125.400 26.200 1185.000 26.800 ;
        RECT 1125.800 25.600 1185.000 26.200 ;
        RECT 1126.200 25.000 1185.000 25.600 ;
        RECT 1126.600 24.400 1185.000 25.000 ;
        RECT 1127.000 23.800 1185.000 24.400 ;
        RECT 1127.400 23.200 1185.000 23.800 ;
        RECT 1127.800 22.600 1185.000 23.200 ;
        RECT 1128.200 22.000 1185.000 22.600 ;
        RECT 1128.600 21.400 1185.000 22.000 ;
        RECT 1129.000 20.800 1185.000 21.400 ;
        RECT 1129.400 20.200 1185.000 20.800 ;
        RECT 1129.800 19.600 1185.000 20.200 ;
        RECT 1130.200 19.000 1185.000 19.600 ;
        RECT 1130.600 18.400 1185.000 19.000 ;
        RECT 1131.000 17.800 1185.000 18.400 ;
        RECT 1131.400 17.200 1185.000 17.800 ;
        RECT 1131.800 16.600 1185.000 17.200 ;
        RECT 1132.200 16.000 1185.000 16.600 ;
        RECT 1132.600 15.400 1185.000 16.000 ;
        RECT 1133.000 14.800 1185.000 15.400 ;
        RECT 1133.400 14.200 1185.000 14.800 ;
        RECT 1133.800 13.600 1185.000 14.200 ;
        RECT 1134.200 13.000 1185.000 13.600 ;
        RECT 1134.600 12.400 1185.000 13.000 ;
  END
END anan_logo
END LIBRARY

